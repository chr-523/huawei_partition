module gated_clk_cell_344 ( clk_in, global_en, module_en, local_en, 
        external_en, pad_yy_icg_scan_en, clk_out );
  input clk_in, global_en, module_en, local_en, external_en,
         pad_yy_icg_scan_en;
  output clk_out;

  wire   clk_in;
  assign clk_out = clk_in;

endmodule


module aq_ifu_pcgen_0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196;

  sky130_fd_sc_hd__inv_1 U2 ( .A(A[20]), .Y(n159) );
  sky130_fd_sc_hd__inv_1 U3 ( .A(A[18]), .Y(n172) );
  sky130_fd_sc_hd__and2_1 U4 ( .A(n102), .B(A[46]), .X(n1) );
  sky130_fd_sc_hd__nand2_2 U5 ( .A(n130), .B(n131), .Y(n91) );
  sky130_fd_sc_hd__inv_2 U6 ( .A(n91), .Y(n112) );
  sky130_fd_sc_hd__nand3_1 U7 ( .A(A[32]), .B(A[33]), .C(n124), .Y(n97) );
  sky130_fd_sc_hd__inv_1 U8 ( .A(A[2]), .Y(SUM[2]) );
  sky130_fd_sc_hd__inv_1 U9 ( .A(A[16]), .Y(n181) );
  sky130_fd_sc_hd__and2_1 U10 ( .A(n70), .B(A[53]), .X(n2) );
  sky130_fd_sc_hd__inv_1 U11 ( .A(A[15]), .Y(n180) );
  sky130_fd_sc_hd__inv_1 U12 ( .A(A[3]), .Y(n196) );
  sky130_fd_sc_hd__nand3_1 U13 ( .A(n160), .B(n161), .C(n162), .Y(n3) );
  sky130_fd_sc_hd__clkinv_1 U14 ( .A(A[28]), .Y(n143) );
  sky130_fd_sc_hd__clkinv_1 U15 ( .A(n67), .Y(n65) );
  sky130_fd_sc_hd__clkinv_1 U16 ( .A(A[31]), .Y(n140) );
  sky130_fd_sc_hd__inv_1 U17 ( .A(n158), .Y(n163) );
  sky130_fd_sc_hd__inv_1 U18 ( .A(n36), .Y(n191) );
  sky130_fd_sc_hd__and2_1 U19 ( .A(A[9]), .B(n35), .X(n22) );
  sky130_fd_sc_hd__and2_1 U20 ( .A(n168), .B(A[20]), .X(n17) );
  sky130_fd_sc_hd__and2_1 U21 ( .A(n22), .B(A[10]), .X(n32) );
  sky130_fd_sc_hd__and2_1 U22 ( .A(A[22]), .B(n14), .X(n164) );
  sky130_fd_sc_hd__clkinv_1 U23 ( .A(n71), .Y(n70) );
  sky130_fd_sc_hd__inv_1 U24 ( .A(n85), .Y(n81) );
  sky130_fd_sc_hd__inv_1 U25 ( .A(n104), .Y(n105) );
  sky130_fd_sc_hd__or2_2 U26 ( .A(n97), .B(n98), .X(n113) );
  sky130_fd_sc_hd__inv_1 U27 ( .A(n91), .Y(n51) );
  sky130_fd_sc_hd__or2_2 U28 ( .A(n97), .B(n91), .X(n6) );
  sky130_fd_sc_hd__or2_2 U29 ( .A(n113), .B(n91), .X(n7) );
  sky130_fd_sc_hd__inv_1 U30 ( .A(n74), .Y(n77) );
  sky130_fd_sc_hd__inv_1 U31 ( .A(n137), .Y(n160) );
  sky130_fd_sc_hd__inv_1 U32 ( .A(n100), .Y(n102) );
  sky130_fd_sc_hd__inv_1 U33 ( .A(A[39]), .Y(n118) );
  sky130_fd_sc_hd__and2_1 U34 ( .A(n171), .B(A[17]), .X(n24) );
  sky130_fd_sc_hd__and2_1 U35 ( .A(n112), .B(A[32]), .X(n13) );
  sky130_fd_sc_hd__and2_1 U36 ( .A(n26), .B(A[5]), .X(n27) );
  sky130_fd_sc_hd__and2_1 U37 ( .A(A[4]), .B(n12), .X(n26) );
  sky130_fd_sc_hd__and2_1 U38 ( .A(A[33]), .B(n13), .X(n126) );
  sky130_fd_sc_hd__and2_1 U39 ( .A(n120), .B(A[37]), .X(n16) );
  sky130_fd_sc_hd__and2_1 U40 ( .A(n5), .B(A[54]), .X(n20) );
  sky130_fd_sc_hd__and2_1 U41 ( .A(n126), .B(A[34]), .X(n19) );
  sky130_fd_sc_hd__and2_1 U42 ( .A(n27), .B(A[6]), .X(n33) );
  sky130_fd_sc_hd__and2_1 U43 ( .A(n16), .B(A[38]), .X(n9) );
  sky130_fd_sc_hd__and2_1 U44 ( .A(n18), .B(A[42]), .X(n21) );
  sky130_fd_sc_hd__and2_1 U45 ( .A(A[18]), .B(n24), .X(n31) );
  sky130_fd_sc_hd__and2_1 U46 ( .A(n4), .B(A[40]), .X(n30) );
  sky130_fd_sc_hd__and2_1 U47 ( .A(n105), .B(A[44]), .X(n8) );
  sky130_fd_sc_hd__and2_1 U48 ( .A(n57), .B(n58), .X(n23) );
  sky130_fd_sc_hd__clkinv_1 U49 ( .A(A[30]), .Y(n141) );
  sky130_fd_sc_hd__clkinv_1 U50 ( .A(A[29]), .Y(n142) );
  sky130_fd_sc_hd__inv_1 U51 ( .A(n38), .Y(n37) );
  sky130_fd_sc_hd__inv_1 U52 ( .A(A[44]), .Y(n106) );
  sky130_fd_sc_hd__inv_1 U53 ( .A(A[45]), .Y(n103) );
  sky130_fd_sc_hd__inv_1 U54 ( .A(A[46]), .Y(n101) );
  sky130_fd_sc_hd__inv_1 U55 ( .A(A[42]), .Y(n110) );
  sky130_fd_sc_hd__inv_1 U56 ( .A(A[6]), .Y(n41) );
  sky130_fd_sc_hd__inv_1 U57 ( .A(A[9]), .Y(n34) );
  sky130_fd_sc_hd__inv_1 U58 ( .A(A[5]), .Y(n54) );
  sky130_fd_sc_hd__inv_1 U59 ( .A(A[4]), .Y(n87) );
  sky130_fd_sc_hd__inv_1 U60 ( .A(A[10]), .Y(n193) );
  sky130_fd_sc_hd__inv_1 U61 ( .A(n179), .Y(n187) );
  sky130_fd_sc_hd__inv_1 U62 ( .A(A[12]), .Y(n190) );
  sky130_fd_sc_hd__inv_1 U63 ( .A(A[41]), .Y(n111) );
  sky130_fd_sc_hd__inv_1 U64 ( .A(A[47]), .Y(n99) );
  sky130_fd_sc_hd__inv_1 U65 ( .A(A[43]), .Y(n109) );
  sky130_fd_sc_hd__inv_1 U66 ( .A(A[11]), .Y(n192) );
  sky130_fd_sc_hd__inv_1 U67 ( .A(n40), .Y(n39) );
  sky130_fd_sc_hd__inv_1 U68 ( .A(A[26]), .Y(n154) );
  sky130_fd_sc_hd__inv_1 U69 ( .A(n115), .Y(n114) );
  sky130_fd_sc_hd__inv_1 U70 ( .A(A[40]), .Y(n115) );
  sky130_fd_sc_hd__inv_1 U71 ( .A(A[50]), .Y(n85) );
  sky130_fd_sc_hd__clkinv_1 U72 ( .A(n116), .Y(n117) );
  sky130_fd_sc_hd__inv_1 U73 ( .A(A[36]), .Y(n116) );
  sky130_fd_sc_hd__inv_1 U74 ( .A(A[56]), .Y(n67) );
  sky130_fd_sc_hd__inv_1 U75 ( .A(n60), .Y(n58) );
  sky130_fd_sc_hd__inv_1 U76 ( .A(n56), .Y(n53) );
  sky130_fd_sc_hd__inv_1 U77 ( .A(A[57]), .Y(n64) );
  sky130_fd_sc_hd__inv_1 U78 ( .A(n150), .Y(n149) );
  sky130_fd_sc_hd__inv_1 U79 ( .A(n162), .Y(n169) );
  sky130_fd_sc_hd__and2_1 U80 ( .A(A[2]), .B(A[3]), .X(n12) );
  sky130_fd_sc_hd__and2_1 U81 ( .A(n147), .B(A[29]), .X(n15) );
  sky130_fd_sc_hd__and2_1 U82 ( .A(A[25]), .B(n155), .X(n153) );
  sky130_fd_sc_hd__and2_1 U83 ( .A(n189), .B(A[12]), .X(n25) );
  sky130_fd_sc_hd__nor2b_1 U84 ( .B_N(A[14]), .A(n176), .Y(n175) );
  sky130_fd_sc_hd__clkinv_1 U85 ( .A(n195), .Y(n40) );
  sky130_fd_sc_hd__inv_1 U86 ( .A(A[7]), .Y(n195) );
  sky130_fd_sc_hd__clkinv_1 U87 ( .A(n194), .Y(n38) );
  sky130_fd_sc_hd__inv_1 U88 ( .A(A[8]), .Y(n194) );
  sky130_fd_sc_hd__clkinv_1 U89 ( .A(n188), .Y(n179) );
  sky130_fd_sc_hd__inv_1 U90 ( .A(A[13]), .Y(n188) );
  sky130_fd_sc_hd__and2_0 U91 ( .A(n112), .B(n107), .X(n4) );
  sky130_fd_sc_hd__inv_2 U92 ( .A(n113), .Y(n107) );
  sky130_fd_sc_hd__nor2_1 U93 ( .A(n3), .B(n144), .Y(n150) );
  sky130_fd_sc_hd__nor2_1 U94 ( .A(n169), .B(n137), .Y(n168) );
  sky130_fd_sc_hd__nor2_1 U95 ( .A(n143), .B(n149), .Y(n147) );
  sky130_fd_sc_hd__nand3_1 U96 ( .A(n107), .B(n108), .C(n112), .Y(n104) );
  sky130_fd_sc_hd__inv_1 U97 ( .A(n93), .Y(n108) );
  sky130_fd_sc_hd__nor2b_1 U98 ( .B_N(n2), .A(n49), .Y(n5) );
  sky130_fd_sc_hd__nor2_1 U99 ( .A(n136), .B(n137), .Y(n135) );
  sky130_fd_sc_hd__nor2_1 U100 ( .A(n142), .B(n143), .Y(n138) );
  sky130_fd_sc_hd__nor2_1 U101 ( .A(n140), .B(n141), .Y(n139) );
  sky130_fd_sc_hd__nand2b_1 U102 ( .A_N(n61), .B(n5), .Y(n62) );
  sky130_fd_sc_hd__inv_2 U103 ( .A(n12), .Y(n132) );
  sky130_fd_sc_hd__inv_1 U104 ( .A(n98), .Y(n95) );
  sky130_fd_sc_hd__inv_1 U105 ( .A(n122), .Y(n120) );
  sky130_fd_sc_hd__nor2_1 U106 ( .A(n116), .B(n97), .Y(n123) );
  sky130_fd_sc_hd__inv_1 U107 ( .A(n145), .Y(n161) );
  sky130_fd_sc_hd__nor2_1 U108 ( .A(n132), .B(n176), .Y(n36) );
  sky130_fd_sc_hd__nor2_1 U109 ( .A(n191), .B(n177), .Y(n189) );
  sky130_fd_sc_hd__nor2_1 U110 ( .A(n90), .B(n71), .Y(n72) );
  sky130_fd_sc_hd__nor2_1 U111 ( .A(n86), .B(n82), .Y(n83) );
  sky130_fd_sc_hd__nor2_1 U112 ( .A(n86), .B(n78), .Y(n79) );
  sky130_fd_sc_hd__nor2_1 U113 ( .A(n86), .B(n77), .Y(n75) );
  sky130_fd_sc_hd__inv_1 U114 ( .A(n97), .Y(n96) );
  sky130_fd_sc_hd__nor2_1 U115 ( .A(n132), .B(n133), .Y(n131) );
  sky130_fd_sc_hd__nor2_1 U116 ( .A(n144), .B(n145), .Y(n134) );
  sky130_fd_sc_hd__nor2_1 U117 ( .A(n132), .B(n133), .Y(n162) );
  sky130_fd_sc_hd__nor2b_1 U118 ( .B_N(A[24]), .A(n3), .Y(n155) );
  sky130_fd_sc_hd__nand3_1 U119 ( .A(A[45]), .B(A[44]), .C(n105), .Y(n100) );
  sky130_fd_sc_hd__nor2_1 U120 ( .A(n49), .B(n11), .Y(n10) );
  sky130_fd_sc_hd__or2_0 U121 ( .A(n47), .B(n48), .X(n11) );
  sky130_fd_sc_hd__and2_0 U122 ( .A(n17), .B(n163), .X(n14) );
  sky130_fd_sc_hd__and3_1 U123 ( .A(A[41]), .B(A[40]), .C(n4), .X(n18) );
  sky130_fd_sc_hd__nor2b_1 U124 ( .B_N(A[51]), .A(n78), .Y(n74) );
  sky130_fd_sc_hd__nor2_1 U125 ( .A(n191), .B(n37), .Y(n35) );
  sky130_fd_sc_hd__nor2b_1 U126 ( .B_N(A[16]), .A(n169), .Y(n171) );
  sky130_fd_sc_hd__nand2b_1 U127 ( .A_N(n82), .B(n81), .Y(n78) );
  sky130_fd_sc_hd__nor2_1 U128 ( .A(n64), .B(n61), .Y(n57) );
  sky130_fd_sc_hd__nor2b_1 U129 ( .B_N(A[48]), .A(n90), .Y(n88) );
  sky130_fd_sc_hd__and2_0 U130 ( .A(A[54]), .B(A[55]), .X(n28) );
  sky130_fd_sc_hd__and2_0 U131 ( .A(n23), .B(n53), .X(n29) );
  sky130_fd_sc_hd__inv_2 U132 ( .A(A[33]), .Y(n128) );
  sky130_fd_sc_hd__and2_0 U133 ( .A(A[35]), .B(A[34]), .X(n124) );
  sky130_fd_sc_hd__inv_2 U134 ( .A(A[22]), .Y(n166) );
  sky130_fd_sc_hd__inv_2 U135 ( .A(A[25]), .Y(n156) );
  sky130_fd_sc_hd__inv_2 U136 ( .A(A[34]), .Y(n127) );
  sky130_fd_sc_hd__inv_2 U137 ( .A(A[24]), .Y(n157) );
  sky130_fd_sc_hd__inv_2 U138 ( .A(A[32]), .Y(n129) );
  sky130_fd_sc_hd__and2_0 U139 ( .A(n179), .B(n25), .X(n184) );
  sky130_fd_sc_hd__inv_2 U140 ( .A(A[51]), .Y(n80) );
  sky130_fd_sc_hd__inv_2 U141 ( .A(A[35]), .Y(n125) );
  sky130_fd_sc_hd__inv_2 U142 ( .A(n163), .Y(n167) );
  sky130_fd_sc_hd__inv_2 U143 ( .A(A[38]), .Y(n119) );
  sky130_fd_sc_hd__inv_2 U144 ( .A(A[37]), .Y(n121) );
  sky130_fd_sc_hd__inv_2 U145 ( .A(A[17]), .Y(n173) );
  sky130_fd_sc_hd__inv_2 U146 ( .A(n64), .Y(n63) );
  sky130_fd_sc_hd__inv_2 U147 ( .A(A[19]), .Y(n170) );
  sky130_fd_sc_hd__inv_2 U148 ( .A(A[23]), .Y(n165) );
  sky130_fd_sc_hd__inv_2 U149 ( .A(A[27]), .Y(n151) );
  sky130_fd_sc_hd__inv_2 U150 ( .A(A[54]), .Y(n69) );
  sky130_fd_sc_hd__inv_2 U151 ( .A(A[55]), .Y(n68) );
  sky130_fd_sc_hd__inv_2 U152 ( .A(A[53]), .Y(n73) );
  sky130_fd_sc_hd__inv_2 U153 ( .A(A[52]), .Y(n76) );
  sky130_fd_sc_hd__inv_2 U154 ( .A(n81), .Y(n84) );
  sky130_fd_sc_hd__inv_2 U155 ( .A(A[49]), .Y(n89) );
  sky130_fd_sc_hd__nor2_1 U156 ( .A(n177), .B(n178), .Y(n174) );
  sky130_fd_sc_hd__nor2b_1 U157 ( .B_N(n10), .A(n44), .Y(n42) );
  sky130_fd_sc_hd__clkinv_1 U158 ( .A(A[21]), .Y(n158) );
  sky130_fd_sc_hd__inv_1 U159 ( .A(A[60]), .Y(n47) );
  sky130_fd_sc_hd__clkinv_1 U160 ( .A(A[58]), .Y(n60) );
  sky130_fd_sc_hd__clkinv_1 U161 ( .A(A[59]), .Y(n56) );
  sky130_fd_sc_hd__inv_1 U162 ( .A(n186), .Y(n185) );
  sky130_fd_sc_hd__inv_1 U163 ( .A(A[14]), .Y(n186) );
  sky130_fd_sc_hd__inv_1 U164 ( .A(A[61]), .Y(n46) );
  sky130_fd_sc_hd__clkinv_1 U165 ( .A(A[63]), .Y(n43) );
  sky130_fd_sc_hd__nand2_1 U166 ( .A(A[61]), .B(n10), .Y(n45) );
  sky130_fd_sc_hd__nand2_1 U167 ( .A(n29), .B(n5), .Y(n52) );
  sky130_fd_sc_hd__nand2_1 U168 ( .A(n15), .B(A[30]), .Y(n146) );
  sky130_fd_sc_hd__nand2_1 U169 ( .A(n153), .B(A[26]), .Y(n152) );
  sky130_fd_sc_hd__nand2_1 U170 ( .A(n184), .B(n185), .Y(n182) );
  sky130_fd_sc_hd__nand2_1 U171 ( .A(n23), .B(n5), .Y(n55) );
  sky130_fd_sc_hd__nand2_1 U172 ( .A(n57), .B(n5), .Y(n59) );
  sky130_fd_sc_hd__nand2_1 U173 ( .A(n28), .B(n5), .Y(n66) );
  sky130_fd_sc_hd__nand2_1 U174 ( .A(n50), .B(n51), .Y(n86) );
  sky130_fd_sc_hd__nand2_1 U175 ( .A(n50), .B(n51), .Y(n90) );
  sky130_fd_sc_hd__nand2_1 U176 ( .A(A[62]), .B(A[61]), .Y(n44) );
  sky130_fd_sc_hd__xnor2_1 U177 ( .A(n34), .B(n35), .Y(SUM[9]) );
  sky130_fd_sc_hd__xnor2_1 U178 ( .A(n36), .B(n37), .Y(SUM[8]) );
  sky130_fd_sc_hd__xnor2_1 U179 ( .A(n33), .B(n39), .Y(SUM[7]) );
  sky130_fd_sc_hd__xnor2_1 U180 ( .A(n41), .B(n27), .Y(SUM[6]) );
  sky130_fd_sc_hd__xnor2_1 U181 ( .A(n42), .B(n43), .Y(SUM[63]) );
  sky130_fd_sc_hd__xnor2_1 U182 ( .A(n45), .B(A[62]), .Y(SUM[62]) );
  sky130_fd_sc_hd__xnor2_1 U183 ( .A(n46), .B(n10), .Y(SUM[61]) );
  sky130_fd_sc_hd__nand2_1 U184 ( .A(n2), .B(n29), .Y(n48) );
  sky130_fd_sc_hd__nand2_1 U185 ( .A(n50), .B(n51), .Y(n49) );
  sky130_fd_sc_hd__xnor2_1 U186 ( .A(n52), .B(A[60]), .Y(SUM[60]) );
  sky130_fd_sc_hd__xnor2_1 U187 ( .A(n54), .B(n26), .Y(SUM[5]) );
  sky130_fd_sc_hd__xnor2_1 U188 ( .A(n55), .B(n53), .Y(SUM[59]) );
  sky130_fd_sc_hd__xnor2_1 U189 ( .A(n59), .B(n58), .Y(SUM[58]) );
  sky130_fd_sc_hd__xnor2_1 U190 ( .A(n62), .B(n63), .Y(SUM[57]) );
  sky130_fd_sc_hd__nand2_1 U191 ( .A(n28), .B(n65), .Y(n61) );
  sky130_fd_sc_hd__xnor2_1 U192 ( .A(n66), .B(n65), .Y(SUM[56]) );
  sky130_fd_sc_hd__xnor2_1 U193 ( .A(n20), .B(n68), .Y(SUM[55]) );
  sky130_fd_sc_hd__xnor2_1 U194 ( .A(n5), .B(n69), .Y(SUM[54]) );
  sky130_fd_sc_hd__xnor2_1 U195 ( .A(n72), .B(n73), .Y(SUM[53]) );
  sky130_fd_sc_hd__nand2_1 U196 ( .A(n74), .B(A[52]), .Y(n71) );
  sky130_fd_sc_hd__xnor2_1 U197 ( .A(n75), .B(n76), .Y(SUM[52]) );
  sky130_fd_sc_hd__xnor2_1 U198 ( .A(n79), .B(n80), .Y(SUM[51]) );
  sky130_fd_sc_hd__xnor2_1 U199 ( .A(n83), .B(n84), .Y(SUM[50]) );
  sky130_fd_sc_hd__nand2_1 U200 ( .A(A[48]), .B(A[49]), .Y(n82) );
  sky130_fd_sc_hd__xnor2_1 U201 ( .A(n12), .B(n87), .Y(SUM[4]) );
  sky130_fd_sc_hd__xnor2_1 U202 ( .A(n88), .B(n89), .Y(SUM[49]) );
  sky130_fd_sc_hd__xnor2_1 U203 ( .A(n90), .B(A[48]), .Y(SUM[48]) );
  sky130_fd_sc_hd__nor3_2 U204 ( .A(n92), .B(n93), .C(n94), .Y(n50) );
  sky130_fd_sc_hd__nand4_1 U205 ( .A(A[44]), .B(A[45]), .C(A[47]), .D(A[46]), 
        .Y(n94) );
  sky130_fd_sc_hd__nand2_1 U206 ( .A(n95), .B(n96), .Y(n92) );
  sky130_fd_sc_hd__xnor2_1 U207 ( .A(n1), .B(n99), .Y(SUM[47]) );
  sky130_fd_sc_hd__xnor2_1 U208 ( .A(n101), .B(n102), .Y(SUM[46]) );
  sky130_fd_sc_hd__xnor2_1 U209 ( .A(n103), .B(n8), .Y(SUM[45]) );
  sky130_fd_sc_hd__xnor2_1 U210 ( .A(n105), .B(n106), .Y(SUM[44]) );
  sky130_fd_sc_hd__nand4_1 U211 ( .A(A[41]), .B(A[40]), .C(A[42]), .D(A[43]), 
        .Y(n93) );
  sky130_fd_sc_hd__xnor2_1 U212 ( .A(n21), .B(n109), .Y(SUM[43]) );
  sky130_fd_sc_hd__xnor2_1 U213 ( .A(n110), .B(n18), .Y(SUM[42]) );
  sky130_fd_sc_hd__xnor2_1 U214 ( .A(n30), .B(n111), .Y(SUM[41]) );
  sky130_fd_sc_hd__xnor2_1 U215 ( .A(n7), .B(n114), .Y(SUM[40]) );
  sky130_fd_sc_hd__nand4_1 U216 ( .A(A[38]), .B(A[39]), .C(A[37]), .D(n117), 
        .Y(n98) );
  sky130_fd_sc_hd__xnor2_1 U217 ( .A(A[2]), .B(n196), .Y(SUM[3]) );
  sky130_fd_sc_hd__xnor2_1 U218 ( .A(n9), .B(n118), .Y(SUM[39]) );
  sky130_fd_sc_hd__xnor2_1 U219 ( .A(n119), .B(n16), .Y(SUM[38]) );
  sky130_fd_sc_hd__xnor2_1 U220 ( .A(n121), .B(n120), .Y(SUM[37]) );
  sky130_fd_sc_hd__nand2_1 U221 ( .A(n123), .B(n112), .Y(n122) );
  sky130_fd_sc_hd__xnor2_1 U222 ( .A(n6), .B(n117), .Y(SUM[36]) );
  sky130_fd_sc_hd__xnor2_1 U223 ( .A(n19), .B(n125), .Y(SUM[35]) );
  sky130_fd_sc_hd__xnor2_1 U224 ( .A(n127), .B(n126), .Y(SUM[34]) );
  sky130_fd_sc_hd__xnor2_1 U225 ( .A(n13), .B(n128), .Y(SUM[33]) );
  sky130_fd_sc_hd__xnor2_1 U226 ( .A(n51), .B(n129), .Y(SUM[32]) );
  sky130_fd_sc_hd__and2_1 U227 ( .A(n134), .B(n135), .X(n130) );
  sky130_fd_sc_hd__nand2_1 U228 ( .A(n138), .B(n139), .Y(n136) );
  sky130_fd_sc_hd__xor2_1 U229 ( .A(n140), .B(n146), .X(SUM[31]) );
  sky130_fd_sc_hd__xnor2_1 U230 ( .A(n141), .B(n15), .Y(SUM[30]) );
  sky130_fd_sc_hd__xnor2_1 U231 ( .A(n142), .B(n147), .Y(SUM[29]) );
  sky130_fd_sc_hd__xnor2_1 U232 ( .A(n150), .B(n143), .Y(SUM[28]) );
  sky130_fd_sc_hd__nand4_1 U233 ( .A(A[25]), .B(A[24]), .C(A[26]), .D(A[27]), 
        .Y(n144) );
  sky130_fd_sc_hd__xor2_1 U234 ( .A(n151), .B(n152), .X(SUM[27]) );
  sky130_fd_sc_hd__xnor2_1 U235 ( .A(n154), .B(n153), .Y(SUM[26]) );
  sky130_fd_sc_hd__xnor2_1 U236 ( .A(n155), .B(n156), .Y(SUM[25]) );
  sky130_fd_sc_hd__xor2_1 U237 ( .A(n157), .B(n3), .X(SUM[24]) );
  sky130_fd_sc_hd__nand4_1 U238 ( .A(A[20]), .B(n163), .C(A[22]), .D(A[23]), 
        .Y(n145) );
  sky130_fd_sc_hd__xnor2_1 U239 ( .A(n164), .B(n165), .Y(SUM[23]) );
  sky130_fd_sc_hd__xnor2_1 U240 ( .A(n14), .B(n166), .Y(SUM[22]) );
  sky130_fd_sc_hd__xnor2_1 U241 ( .A(n167), .B(n17), .Y(SUM[21]) );
  sky130_fd_sc_hd__xnor2_1 U242 ( .A(n159), .B(n168), .Y(SUM[20]) );
  sky130_fd_sc_hd__nand4_1 U243 ( .A(A[18]), .B(A[19]), .C(A[17]), .D(A[16]), 
        .Y(n137) );
  sky130_fd_sc_hd__xnor2_1 U244 ( .A(n31), .B(n170), .Y(SUM[19]) );
  sky130_fd_sc_hd__xnor2_1 U245 ( .A(n172), .B(n24), .Y(SUM[18]) );
  sky130_fd_sc_hd__xnor2_1 U246 ( .A(n173), .B(n171), .Y(SUM[17]) );
  sky130_fd_sc_hd__xor2_1 U247 ( .A(n181), .B(n169), .X(SUM[16]) );
  sky130_fd_sc_hd__nand2_1 U248 ( .A(n174), .B(n175), .Y(n133) );
  sky130_fd_sc_hd__nand3_1 U249 ( .A(n179), .B(A[12]), .C(A[15]), .Y(n178) );
  sky130_fd_sc_hd__xnor2_1 U250 ( .A(n182), .B(n183), .Y(SUM[15]) );
  sky130_fd_sc_hd__inv_1 U251 ( .A(n180), .Y(n183) );
  sky130_fd_sc_hd__xnor2_1 U252 ( .A(n186), .B(n184), .Y(SUM[14]) );
  sky130_fd_sc_hd__xnor2_1 U253 ( .A(n25), .B(n187), .Y(SUM[13]) );
  sky130_fd_sc_hd__xnor2_1 U254 ( .A(n189), .B(n190), .Y(SUM[12]) );
  sky130_fd_sc_hd__nand4_1 U255 ( .A(A[9]), .B(n38), .C(A[10]), .D(A[11]), .Y(
        n177) );
  sky130_fd_sc_hd__xnor2_1 U256 ( .A(n32), .B(n192), .Y(SUM[11]) );
  sky130_fd_sc_hd__xnor2_1 U257 ( .A(n22), .B(n193), .Y(SUM[10]) );
  sky130_fd_sc_hd__nand4_1 U258 ( .A(A[5]), .B(A[4]), .C(A[6]), .D(n40), .Y(
        n176) );
endmodule


module aq_ifu_pcgen_0 ( btb_pcgen_tar_pc, btb_xx_chgflw_vld, cp0_ifu_icg_en, 
        cp0_xx_mrvbr, cp0_yy_clk_en, cpurst_b, forever_cpuclk, 
        icache_pcgen_addr, icache_pcgen_grant, icache_pcgen_grant_gate, 
        icache_pcgen_inst_vld, icache_pcgen_inst_vld_gate, ifu_iu_chgflw_pc, 
        ifu_iu_chgflw_vld, ipack_pcgen_reissue, iu_ifu_tar_pc, 
        iu_ifu_tar_pc_vld, iu_ifu_tar_pc_vld_gate, pad_yy_icg_scan_en, 
        pcgen_btb_ifpc, pcgen_ctrl_chgflw_vld, pcgen_ibuf_chgflw_vld, 
        pcgen_icache_chgflw_vld, pcgen_icache_seq_tag, pcgen_icache_va, 
        pcgen_pred_flush_vld, pcgen_pred_ifpc, pcgen_top_buf_chgflw, 
        pred_pcgen_chgflw_pc, pred_pcgen_chgflw_vld, 
        pred_pcgen_chgflw_vld_gate, pred_pcgen_curflw_pc, 
        pred_pcgen_curflw_vld, pred_pcgen_curflw_vld_gate, rtu_ifu_chgflw_pc, 
        rtu_ifu_chgflw_vld, vec_pcgen_idle, vec_pcgen_rst_vld );
  input [39:0] btb_pcgen_tar_pc;
  input [39:0] cp0_xx_mrvbr;
  input [39:0] icache_pcgen_addr;
  output [39:0] ifu_iu_chgflw_pc;
  input [63:0] iu_ifu_tar_pc;
  output [39:0] pcgen_btb_ifpc;
  output [33:0] pcgen_icache_seq_tag;
  output [63:0] pcgen_icache_va;
  output [39:0] pcgen_pred_ifpc;
  input [39:0] pred_pcgen_chgflw_pc;
  input [39:0] pred_pcgen_curflw_pc;
  input [39:0] rtu_ifu_chgflw_pc;
  input btb_xx_chgflw_vld, cp0_ifu_icg_en, cp0_yy_clk_en, cpurst_b,
         forever_cpuclk, icache_pcgen_grant, icache_pcgen_grant_gate,
         icache_pcgen_inst_vld, icache_pcgen_inst_vld_gate,
         ipack_pcgen_reissue, iu_ifu_tar_pc_vld, iu_ifu_tar_pc_vld_gate,
         pad_yy_icg_scan_en, pred_pcgen_chgflw_vld, pred_pcgen_chgflw_vld_gate,
         pred_pcgen_curflw_vld, pred_pcgen_curflw_vld_gate, rtu_ifu_chgflw_vld,
         vec_pcgen_idle, vec_pcgen_rst_vld;
  output ifu_iu_chgflw_vld, pcgen_ctrl_chgflw_vld, pcgen_ibuf_chgflw_vld,
         pcgen_icache_chgflw_vld, pcgen_pred_flush_vld, pcgen_top_buf_chgflw;
  wire   n_Logic1_, n1, pcgen_icg_en, pcgen_ifpc_5, pcgen_ifpc_4, pcgen_ifpc_3,
         pcgen_ifpc_2, pcgen_ifpc_1, pcgen_ifpc_0, N22, N23, N24, N25, N26,
         N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54,
         N55, N56, N57, N58, N59, N60, N61, N85, N86, N87, N88, N89, N90, N91,
         N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104,
         N105, N106, N107, N108, n180, n181, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, pcgen_pred_flush_vld, n533,
         __UC__n_1, __UC__n_2;
  wire   [63:40] pcgen_ifpc;
  wire   [63:2] pcgen_ifpc_inc;
  wire   forever_cpuclk;
  wire   pcgen_cpuclk;
  assign pcgen_icache_seq_tag[33] = pcgen_btb_ifpc[39];
  assign pcgen_icache_seq_tag[32] = pcgen_btb_ifpc[38];
  assign pcgen_icache_seq_tag[31] = pcgen_btb_ifpc[37];
  assign pcgen_icache_seq_tag[30] = pcgen_btb_ifpc[36];
  assign pcgen_icache_seq_tag[29] = pcgen_btb_ifpc[35];
  assign pcgen_icache_seq_tag[28] = pcgen_btb_ifpc[34];
  assign pcgen_icache_seq_tag[27] = pcgen_btb_ifpc[33];
  assign pcgen_icache_seq_tag[26] = pcgen_btb_ifpc[32];
  assign pcgen_icache_seq_tag[25] = pcgen_btb_ifpc[31];
  assign pcgen_icache_seq_tag[24] = pcgen_btb_ifpc[30];
  assign pcgen_icache_seq_tag[23] = pcgen_btb_ifpc[29];
  assign pcgen_icache_seq_tag[22] = pcgen_btb_ifpc[28];
  assign pcgen_icache_seq_tag[21] = pcgen_btb_ifpc[27];
  assign pcgen_icache_seq_tag[20] = pcgen_btb_ifpc[26];
  assign pcgen_icache_seq_tag[19] = pcgen_btb_ifpc[25];
  assign pcgen_icache_seq_tag[18] = pcgen_btb_ifpc[24];
  assign pcgen_icache_seq_tag[17] = pcgen_btb_ifpc[23];
  assign pcgen_icache_seq_tag[16] = pcgen_btb_ifpc[22];
  assign pcgen_icache_seq_tag[15] = pcgen_btb_ifpc[21];
  assign pcgen_icache_seq_tag[14] = pcgen_btb_ifpc[20];
  assign pcgen_icache_seq_tag[13] = pcgen_btb_ifpc[19];
  assign pcgen_icache_seq_tag[12] = pcgen_btb_ifpc[18];
  assign pcgen_icache_seq_tag[11] = pcgen_btb_ifpc[17];
  assign pcgen_icache_seq_tag[10] = pcgen_btb_ifpc[16];
  assign pcgen_icache_va[15] = pcgen_btb_ifpc[15];
  assign pcgen_icache_va[14] = pcgen_btb_ifpc[14];
  assign pcgen_icache_va[13] = pcgen_btb_ifpc[13];
  assign pcgen_icache_va[12] = pcgen_btb_ifpc[12];
  assign pcgen_icache_va[11] = pcgen_btb_ifpc[11];
  assign pcgen_icache_va[10] = pcgen_btb_ifpc[10];
  assign pcgen_icache_va[9] = pcgen_btb_ifpc[9];
  assign pcgen_icache_va[8] = pcgen_btb_ifpc[8];
  assign pcgen_icache_va[7] = pcgen_btb_ifpc[7];
  assign pcgen_icache_va[6] = pcgen_btb_ifpc[6];
  assign pcgen_icache_va[5] = pcgen_btb_ifpc[5];
  assign pcgen_icache_va[4] = pcgen_btb_ifpc[4];
  assign pcgen_icache_va[3] = pcgen_btb_ifpc[3];
  assign pcgen_icache_va[2] = pcgen_btb_ifpc[2];
  assign pcgen_icache_va[1] = pcgen_btb_ifpc[1];
  assign pcgen_icache_va[0] = pcgen_btb_ifpc[0];
  assign pcgen_ibuf_chgflw_vld = pcgen_pred_flush_vld;

  sky130_fd_sc_hd__dfrtp_1 pcgen_buf_chgflw_reg ( .D(n533), .CLK(pcgen_cpuclk), 
        .RESET_B(cpurst_b), .Q(pcgen_top_buf_chgflw) );
  gated_clk_cell_344 x_ifu_pcgen_icg_cell ( .clk_in(forever_cpuclk), 
        .global_en(cp0_yy_clk_en), .module_en(cp0_ifu_icg_en), .local_en(
        pcgen_icg_en), .external_en(n1), .pad_yy_icg_scan_en(
        pad_yy_icg_scan_en), .clk_out(pcgen_cpuclk) );
  aq_ifu_pcgen_0_DW01_add_1 add_277 ( .A({pcgen_icache_va[63:16], 
        pcgen_btb_ifpc[15:2], n1, n1}), .B({n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n_Logic1_, n1, n1}), .CI(n1), .SUM({pcgen_ifpc_inc, 
        __UC__n_1, __UC__n_2}) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_0_ ( .D(n433), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[0]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_39_ ( .D(n472), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[39]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_1_ ( .D(n434), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[1]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_38_ ( .D(n471), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[38]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_37_ ( .D(n470), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[37]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_36_ ( .D(n469), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[36]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_35_ ( .D(n468), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[35]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_34_ ( .D(n467), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[34]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_33_ ( .D(n466), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[33]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_32_ ( .D(n465), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[32]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_31_ ( .D(n464), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[31]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_30_ ( .D(n463), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[30]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_29_ ( .D(n462), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[29]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_28_ ( .D(n461), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[28]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_27_ ( .D(n460), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[27]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_26_ ( .D(n459), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[26]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_25_ ( .D(n458), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[25]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_24_ ( .D(n457), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[24]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_23_ ( .D(n456), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[23]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_22_ ( .D(n455), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[22]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_21_ ( .D(n454), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[21]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_20_ ( .D(n453), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[20]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_19_ ( .D(n452), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[19]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_18_ ( .D(n451), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[18]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_17_ ( .D(n450), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[17]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_16_ ( .D(n449), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[16]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_61_ ( .D(N106), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[61]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_62_ ( .D(N107), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[62]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_63_ ( .D(N108), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[63]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_58_ ( .D(N103), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[58]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_52_ ( .D(N97), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[52]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_60_ ( .D(N105), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[60]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_57_ ( .D(N102), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[57]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_59_ ( .D(N104), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[59]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_56_ ( .D(N101), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[56]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_53_ ( .D(N98), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[53]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_51_ ( .D(N96), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[51]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_47_ ( .D(N92), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[47]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_50_ ( .D(N95), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[50]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_55_ ( .D(N100), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[55]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_45_ ( .D(N90), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[45]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_46_ ( .D(N91), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[46]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_43_ ( .D(N88), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[43]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_44_ ( .D(N89), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[44]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_54_ ( .D(N99), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[54]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_49_ ( .D(N94), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[49]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_41_ ( .D(N86), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[41]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_42_ ( .D(N87), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[42]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_48_ ( .D(N93), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[48]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_40_ ( .D(N85), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc[40]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_0_ ( .D(N22), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc_0) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_1_ ( .D(N23), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc_1) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_3_ ( .D(N25), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc_3) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_5_ ( .D(N27), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc_5) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_4_ ( .D(N26), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc_4) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_2_ ( .D(N24), .CLK(pcgen_cpuclk), 
        .Q(pcgen_ifpc_2) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_6_ ( .D(N28), .CLK(pcgen_cpuclk), 
        .Q(pcgen_icache_seq_tag[0]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_14_ ( .D(N36), .CLK(pcgen_cpuclk), 
        .Q(pcgen_icache_seq_tag[8]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_12_ ( .D(N34), .CLK(pcgen_cpuclk), 
        .Q(pcgen_icache_seq_tag[6]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_15_ ( .D(N37), .CLK(pcgen_cpuclk), 
        .Q(pcgen_icache_seq_tag[9]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_13_ ( .D(N35), .CLK(pcgen_cpuclk), 
        .Q(pcgen_icache_seq_tag[7]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_11_ ( .D(N33), .CLK(pcgen_cpuclk), 
        .Q(pcgen_icache_seq_tag[5]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_9_ ( .D(N31), .CLK(pcgen_cpuclk), 
        .Q(pcgen_icache_seq_tag[3]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_10_ ( .D(N32), .CLK(pcgen_cpuclk), 
        .Q(pcgen_icache_seq_tag[4]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_8_ ( .D(N30), .CLK(pcgen_cpuclk), 
        .Q(pcgen_icache_seq_tag[2]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_39_ ( .D(N61), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[39]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_7_ ( .D(N29), .CLK(pcgen_cpuclk), 
        .Q(pcgen_icache_seq_tag[1]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_20_ ( .D(N42), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[20]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_23_ ( .D(N45), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[23]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_27_ ( .D(N49), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[27]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_21_ ( .D(N43), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[21]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_22_ ( .D(N44), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[22]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_18_ ( .D(N40), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[18]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_24_ ( .D(N46), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[24]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_19_ ( .D(N41), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[19]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_16_ ( .D(N38), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[16]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_17_ ( .D(N39), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[17]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_28_ ( .D(N50), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[28]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_30_ ( .D(N52), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[30]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_29_ ( .D(N51), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[29]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_32_ ( .D(N54), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[32]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_38_ ( .D(N60), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[38]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_36_ ( .D(N58), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[36]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_33_ ( .D(N55), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[33]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_37_ ( .D(N59), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[37]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_35_ ( .D(N57), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[35]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_34_ ( .D(N56), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[34]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_25_ ( .D(N47), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[25]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_31_ ( .D(N53), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[31]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_ifpc_reg_26_ ( .D(N48), .CLK(pcgen_cpuclk), 
        .Q(pcgen_btb_ifpc[26]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_14_ ( .D(n447), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[14]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_7_ ( .D(n440), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[7]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_5_ ( .D(n438), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[5]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_12_ ( .D(n445), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[12]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_13_ ( .D(n446), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[13]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_8_ ( .D(n441), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[8]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_9_ ( .D(n442), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[9]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_6_ ( .D(n439), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[6]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_10_ ( .D(n443), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[10]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_11_ ( .D(n444), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[11]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_15_ ( .D(n448), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[15]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_2_ ( .D(n435), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[2]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_4_ ( .D(n437), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[4]) );
  sky130_fd_sc_hd__dfxtp_1 pcgen_pipe_ifpc_reg_3_ ( .D(n436), .CLK(
        pcgen_cpuclk), .Q(pcgen_pred_ifpc[3]) );
  sky130_fd_sc_hd__buf_2 U3 ( .A(n490), .X(n17) );
  sky130_fd_sc_hd__buf_6 U4 ( .A(n366), .X(n85) );
  sky130_fd_sc_hd__buf_2 U5 ( .A(n99), .X(n98) );
  sky130_fd_sc_hd__inv_1 U6 ( .A(vec_pcgen_rst_vld), .Y(n102) );
  sky130_fd_sc_hd__clkbuf_2 U7 ( .A(n103), .X(n97) );
  sky130_fd_sc_hd__dlygate4sd1_1 U8 ( .A(n102), .X(n99) );
  sky130_fd_sc_hd__inv_1 U9 ( .A(ifu_iu_chgflw_vld), .Y(n58) );
  sky130_fd_sc_hd__bufinv_8 U10 ( .A(n106), .Y(ifu_iu_chgflw_vld) );
  sky130_fd_sc_hd__and2_2 U11 ( .A(n25), .B(n100), .X(n2) );
  sky130_fd_sc_hd__buf_2 U12 ( .A(n219), .X(n65) );
  sky130_fd_sc_hd__buf_2 U13 ( .A(n219), .X(n66) );
  sky130_fd_sc_hd__buf_4 U14 ( .A(n219), .X(n64) );
  sky130_fd_sc_hd__and2_4 U15 ( .A(n113), .B(n111), .X(n53) );
  sky130_fd_sc_hd__buf_6 U16 ( .A(n357), .X(n69) );
  sky130_fd_sc_hd__buf_2 U17 ( .A(n51), .X(n79) );
  sky130_fd_sc_hd__buf_1 U18 ( .A(n12), .X(n78) );
  sky130_fd_sc_hd__buf_2 U19 ( .A(n366), .X(n87) );
  sky130_fd_sc_hd__inv_2 U20 ( .A(n85), .Y(n39) );
  sky130_fd_sc_hd__inv_1 U21 ( .A(iu_ifu_tar_pc_vld), .Y(n104) );
  sky130_fd_sc_hd__inv_2 U22 ( .A(n109), .Y(n361) );
  sky130_fd_sc_hd__and2_2 U23 ( .A(iu_ifu_tar_pc_vld), .B(n106), .X(n54) );
  sky130_fd_sc_hd__nand2b_1 U24 ( .A_N(n143), .B(n115), .Y(n139) );
  sky130_fd_sc_hd__and4b_1 U25 ( .B(n104), .C(n106), .D(n488), .A_N(
        pred_pcgen_curflw_vld), .X(n55) );
  sky130_fd_sc_hd__clkinv_1 U26 ( .A(n139), .Y(n120) );
  sky130_fd_sc_hd__a221oi_1 U27 ( .A1(pcgen_ifpc_inc[11]), .A2(n12), .B1(n18), 
        .B2(pcgen_btb_ifpc[11]), .C1(n333), .Y(n3) );
  sky130_fd_sc_hd__inv_2 U28 ( .A(n119), .Y(n115) );
  sky130_fd_sc_hd__a221oi_1 U29 ( .A1(pcgen_ifpc_inc[5]), .A2(n12), .B1(n364), 
        .B2(pcgen_btb_ifpc[5]), .C1(n352), .Y(n4) );
  sky130_fd_sc_hd__a221oi_1 U30 ( .A1(pcgen_ifpc_inc[3]), .A2(n12), .B1(n364), 
        .B2(pcgen_btb_ifpc[3]), .C1(n360), .Y(n5) );
  sky130_fd_sc_hd__a221oi_1 U31 ( .A1(pcgen_ifpc_inc[6]), .A2(n51), .B1(n18), 
        .B2(pcgen_btb_ifpc[6]), .C1(n349), .Y(n6) );
  sky130_fd_sc_hd__mux2_1 U32 ( .A0(n326), .A1(n390), .S(n94), .X(n7) );
  sky130_fd_sc_hd__inv_1 U33 ( .A(vec_pcgen_rst_vld), .Y(n103) );
  sky130_fd_sc_hd__inv_2 U34 ( .A(n88), .Y(n8) );
  sky130_fd_sc_hd__inv_1 U35 ( .A(n11), .Y(n9) );
  sky130_fd_sc_hd__buf_4 U36 ( .A(n479), .X(n88) );
  sky130_fd_sc_hd__clkbuf_2 U37 ( .A(n480), .X(n11) );
  sky130_fd_sc_hd__buf_2 U38 ( .A(n480), .X(n10) );
  sky130_fd_sc_hd__inv_2 U39 ( .A(n486), .Y(n480) );
  sky130_fd_sc_hd__clkbuf_2 U40 ( .A(n361), .X(n72) );
  sky130_fd_sc_hd__and3_4 U41 ( .A(n29), .B(n115), .C(icache_pcgen_grant), .X(
        n12) );
  sky130_fd_sc_hd__nand2_1 U42 ( .A(n87), .B(pcgen_ifpc_5), .Y(n13) );
  sky130_fd_sc_hd__nand2_1 U43 ( .A(icache_pcgen_addr[5]), .B(n84), .Y(n14) );
  sky130_fd_sc_hd__nand3_1 U44 ( .A(n13), .B(n14), .C(n4), .Y(N27) );
  sky130_fd_sc_hd__nand2_1 U45 ( .A(n85), .B(pcgen_ifpc_3), .Y(n15) );
  sky130_fd_sc_hd__nand2_1 U46 ( .A(icache_pcgen_addr[3]), .B(n84), .Y(n16) );
  sky130_fd_sc_hd__nand3_1 U47 ( .A(n15), .B(n16), .C(n5), .Y(N25) );
  sky130_fd_sc_hd__nand2_4 U48 ( .A(n117), .B(n118), .Y(n18) );
  sky130_fd_sc_hd__nand2_4 U49 ( .A(n117), .B(n118), .Y(n364) );
  sky130_fd_sc_hd__nand2_1 U50 ( .A(n86), .B(pcgen_icache_seq_tag[5]), .Y(n19)
         );
  sky130_fd_sc_hd__nand2_1 U51 ( .A(icache_pcgen_addr[11]), .B(n84), .Y(n20)
         );
  sky130_fd_sc_hd__nand3_1 U52 ( .A(n19), .B(n20), .C(n3), .Y(N33) );
  sky130_fd_sc_hd__nand2_1 U53 ( .A(n52), .B(n113), .Y(n21) );
  sky130_fd_sc_hd__nand3_2 U54 ( .A(n143), .B(n124), .C(n22), .Y(n118) );
  sky130_fd_sc_hd__inv_2 U55 ( .A(n21), .Y(n22) );
  sky130_fd_sc_hd__buf_6 U56 ( .A(n49), .X(n84) );
  sky130_fd_sc_hd__inv_1 U57 ( .A(n112), .Y(n113) );
  sky130_fd_sc_hd__nand2_1 U58 ( .A(n490), .B(n55), .Y(pcgen_ctrl_chgflw_vld)
         );
  sky130_fd_sc_hd__nand2_1 U59 ( .A(pcgen_ifpc_inc[13]), .B(n79), .Y(n23) );
  sky130_fd_sc_hd__nand2_1 U60 ( .A(n18), .B(pcgen_btb_ifpc[13]), .Y(n24) );
  sky130_fd_sc_hd__nand3_1 U61 ( .A(n23), .B(n24), .C(n7), .Y(n327) );
  sky130_fd_sc_hd__buf_2 U62 ( .A(n54), .X(n25) );
  sky130_fd_sc_hd__buf_2 U63 ( .A(n54), .X(n26) );
  sky130_fd_sc_hd__buf_2 U64 ( .A(n54), .X(n77) );
  sky130_fd_sc_hd__buf_2 U65 ( .A(n479), .X(n27) );
  sky130_fd_sc_hd__inv_1 U66 ( .A(n485), .Y(n479) );
  sky130_fd_sc_hd__buf_2 U67 ( .A(n361), .X(n71) );
  sky130_fd_sc_hd__buf_2 U68 ( .A(n361), .X(n74) );
  sky130_fd_sc_hd__buf_2 U69 ( .A(n479), .X(n89) );
  sky130_fd_sc_hd__buf_2 U70 ( .A(n479), .X(n90) );
  sky130_fd_sc_hd__inv_1 U71 ( .A(pcgen_icache_seq_tag[3]), .Y(n40) );
  sky130_fd_sc_hd__inv_1 U72 ( .A(pcgen_icache_seq_tag[4]), .Y(n36) );
  sky130_fd_sc_hd__inv_1 U73 ( .A(pcgen_icache_seq_tag[2]), .Y(n33) );
  sky130_fd_sc_hd__inv_1 U74 ( .A(icache_pcgen_addr[8]), .Y(n34) );
  sky130_fd_sc_hd__inv_1 U75 ( .A(icache_pcgen_addr[9]), .Y(n41) );
  sky130_fd_sc_hd__inv_1 U76 ( .A(icache_pcgen_addr[10]), .Y(n37) );
  sky130_fd_sc_hd__buf_6 U77 ( .A(n361), .X(n73) );
  sky130_fd_sc_hd__inv_1 U78 ( .A(n31), .Y(n28) );
  sky130_fd_sc_hd__clkinv_1 U79 ( .A(pred_pcgen_chgflw_vld), .Y(n490) );
  sky130_fd_sc_hd__and2_2 U80 ( .A(n117), .B(n118), .X(n30) );
  sky130_fd_sc_hd__nand2_1 U81 ( .A(ipack_pcgen_reissue), .B(
        icache_pcgen_inst_vld), .Y(n29) );
  sky130_fd_sc_hd__nand2_1 U82 ( .A(ipack_pcgen_reissue), .B(
        icache_pcgen_inst_vld), .Y(n143) );
  sky130_fd_sc_hd__inv_2 U83 ( .A(icache_pcgen_grant), .Y(n124) );
  sky130_fd_sc_hd__buf_6 U84 ( .A(n366), .X(n86) );
  sky130_fd_sc_hd__nand2_2 U85 ( .A(n69), .B(n124), .Y(n137) );
  sky130_fd_sc_hd__inv_1 U86 ( .A(n17), .Y(n31) );
  sky130_fd_sc_hd__dlymetal6s2s_1 U87 ( .A(n12), .X(n32) );
  sky130_fd_sc_hd__dlymetal6s2s_1 U88 ( .A(n12), .X(n80) );
  sky130_fd_sc_hd__dlymetal6s2s_1 U89 ( .A(n51), .X(n81) );
  sky130_fd_sc_hd__o221ai_2 U90 ( .A1(n39), .A2(n33), .B1(n34), .B2(n42), .C1(
        n35), .Y(N30) );
  sky130_fd_sc_hd__a221oi_1 U91 ( .A1(pcgen_ifpc_inc[8]), .A2(n51), .B1(n18), 
        .B2(pcgen_btb_ifpc[8]), .C1(n342), .Y(n35) );
  sky130_fd_sc_hd__bufinv_16 U92 ( .A(n84), .Y(n42) );
  sky130_fd_sc_hd__o221ai_1 U93 ( .A1(n39), .A2(n36), .B1(n37), .B2(n42), .C1(
        n38), .Y(N32) );
  sky130_fd_sc_hd__a221oi_1 U94 ( .A1(pcgen_ifpc_inc[10]), .A2(n12), .B1(n18), 
        .B2(pcgen_btb_ifpc[10]), .C1(n336), .Y(n38) );
  sky130_fd_sc_hd__o221ai_1 U95 ( .A1(n39), .A2(n40), .B1(n41), .B2(n42), .C1(
        n43), .Y(N31) );
  sky130_fd_sc_hd__a221oi_1 U96 ( .A1(pcgen_ifpc_inc[9]), .A2(n51), .B1(n18), 
        .B2(pcgen_btb_ifpc[9]), .C1(n339), .Y(n43) );
  sky130_fd_sc_hd__nand2_1 U97 ( .A(n87), .B(pcgen_icache_seq_tag[6]), .Y(n44)
         );
  sky130_fd_sc_hd__nand2_1 U98 ( .A(icache_pcgen_addr[12]), .B(n84), .Y(n45)
         );
  sky130_fd_sc_hd__nand3_1 U99 ( .A(n44), .B(n45), .C(n46), .Y(N34) );
  sky130_fd_sc_hd__a221oi_1 U100 ( .A1(pcgen_ifpc_inc[12]), .A2(n79), .B1(n18), 
        .B2(pcgen_btb_ifpc[12]), .C1(n330), .Y(n46) );
  sky130_fd_sc_hd__nand2_1 U101 ( .A(n85), .B(pcgen_icache_seq_tag[0]), .Y(n47) );
  sky130_fd_sc_hd__nand2_1 U102 ( .A(icache_pcgen_addr[6]), .B(n84), .Y(n48)
         );
  sky130_fd_sc_hd__nand3_1 U103 ( .A(n47), .B(n48), .C(n6), .Y(N28) );
  sky130_fd_sc_hd__nand2_4 U104 ( .A(n116), .B(n115), .Y(n117) );
  sky130_fd_sc_hd__and3_4 U105 ( .A(n29), .B(n115), .C(icache_pcgen_grant), 
        .X(n51) );
  sky130_fd_sc_hd__inv_1 U106 ( .A(n216), .Y(n61) );
  sky130_fd_sc_hd__inv_1 U107 ( .A(n58), .Y(n57) );
  sky130_fd_sc_hd__inv_1 U108 ( .A(n111), .Y(n357) );
  sky130_fd_sc_hd__clkbuf_1 U109 ( .A(n102), .X(n100) );
  sky130_fd_sc_hd__and2_1 U110 ( .A(pred_pcgen_chgflw_pc[39]), .B(n73), .X(n50) );
  sky130_fd_sc_hd__and2_1 U111 ( .A(n120), .B(n137), .X(n49) );
  sky130_fd_sc_hd__clkbuf_1 U112 ( .A(n102), .X(n101) );
  sky130_fd_sc_hd__and2_1 U113 ( .A(rtu_ifu_chgflw_pc[39]), .B(
        ifu_iu_chgflw_vld), .X(n56) );
  sky130_fd_sc_hd__buf_2 U114 ( .A(n480), .X(n92) );
  sky130_fd_sc_hd__buf_2 U115 ( .A(n480), .X(n93) );
  sky130_fd_sc_hd__buf_2 U116 ( .A(n480), .X(n91) );
  sky130_fd_sc_hd__buf_2 U117 ( .A(n49), .X(n83) );
  sky130_fd_sc_hd__buf_2 U118 ( .A(n49), .X(n82) );
  sky130_fd_sc_hd__inv_1 U119 ( .A(n533), .Y(n114) );
  sky130_fd_sc_hd__inv_2 U120 ( .A(pcgen_pred_flush_vld), .Y(n108) );
  sky130_fd_sc_hd__buf_2 U121 ( .A(n53), .X(n67) );
  sky130_fd_sc_hd__buf_2 U122 ( .A(n54), .X(n75) );
  sky130_fd_sc_hd__buf_2 U123 ( .A(n53), .X(n68) );
  sky130_fd_sc_hd__buf_2 U124 ( .A(n54), .X(n76) );
  sky130_fd_sc_hd__buf_1 U125 ( .A(n357), .X(n70) );
  sky130_fd_sc_hd__inv_2 U126 ( .A(n64), .Y(n63) );
  sky130_fd_sc_hd__inv_2 U127 ( .A(n64), .Y(n62) );
  sky130_fd_sc_hd__inv_2 U128 ( .A(n97), .Y(n94) );
  sky130_fd_sc_hd__and3_1 U129 ( .A(n111), .B(n102), .C(n114), .X(n52) );
  sky130_fd_sc_hd__inv_2 U130 ( .A(n223), .Y(n366) );
  sky130_fd_sc_hd__inv_2 U131 ( .A(n61), .Y(n59) );
  sky130_fd_sc_hd__inv_2 U132 ( .A(n61), .Y(n60) );
  sky130_fd_sc_hd__inv_2 U133 ( .A(n97), .Y(n95) );
  sky130_fd_sc_hd__inv_2 U134 ( .A(n97), .Y(n96) );
  sky130_fd_sc_hd__inv_2 U135 ( .A(rtu_ifu_chgflw_vld), .Y(n106) );
  sky130_fd_sc_hd__inv_1 U136 ( .A(n483), .Y(n220) );
  sky130_fd_sc_hd__nor3_1 U137 ( .A(pred_pcgen_chgflw_vld_gate), .B(n96), .C(
        pred_pcgen_curflw_vld_gate), .Y(n180) );
  sky130_fd_sc_hd__inv_1 U138 ( .A(pcgen_icache_va[63]), .Y(n145) );
  sky130_fd_sc_hd__inv_1 U139 ( .A(pcgen_icache_va[62]), .Y(n148) );
  sky130_fd_sc_hd__inv_1 U140 ( .A(pcgen_icache_va[61]), .Y(n151) );
  sky130_fd_sc_hd__inv_1 U141 ( .A(pcgen_icache_va[60]), .Y(n154) );
  sky130_fd_sc_hd__inv_1 U142 ( .A(pcgen_icache_va[59]), .Y(n157) );
  sky130_fd_sc_hd__inv_1 U143 ( .A(pcgen_icache_va[58]), .Y(n160) );
  sky130_fd_sc_hd__inv_1 U144 ( .A(pcgen_icache_va[55]), .Y(n169) );
  sky130_fd_sc_hd__inv_1 U145 ( .A(pcgen_icache_va[54]), .Y(n172) );
  sky130_fd_sc_hd__inv_1 U146 ( .A(pcgen_icache_va[53]), .Y(n175) );
  sky130_fd_sc_hd__inv_1 U147 ( .A(pcgen_icache_va[52]), .Y(n178) );
  sky130_fd_sc_hd__inv_1 U148 ( .A(pcgen_icache_va[51]), .Y(n183) );
  sky130_fd_sc_hd__inv_1 U149 ( .A(pcgen_icache_va[50]), .Y(n186) );
  sky130_fd_sc_hd__inv_1 U150 ( .A(pcgen_icache_va[49]), .Y(n189) );
  sky130_fd_sc_hd__inv_1 U151 ( .A(pcgen_icache_va[48]), .Y(n192) );
  sky130_fd_sc_hd__inv_1 U152 ( .A(pcgen_icache_va[47]), .Y(n195) );
  sky130_fd_sc_hd__inv_1 U153 ( .A(pcgen_icache_va[46]), .Y(n198) );
  sky130_fd_sc_hd__inv_1 U154 ( .A(pcgen_icache_va[45]), .Y(n201) );
  sky130_fd_sc_hd__inv_1 U155 ( .A(pcgen_icache_va[44]), .Y(n204) );
  sky130_fd_sc_hd__inv_1 U156 ( .A(pcgen_icache_va[43]), .Y(n207) );
  sky130_fd_sc_hd__inv_1 U157 ( .A(pcgen_icache_va[42]), .Y(n210) );
  sky130_fd_sc_hd__inv_1 U158 ( .A(pcgen_icache_va[41]), .Y(n213) );
  sky130_fd_sc_hd__inv_1 U159 ( .A(pcgen_icache_va[40]), .Y(n217) );
  sky130_fd_sc_hd__inv_1 U160 ( .A(pcgen_icache_va[57]), .Y(n163) );
  sky130_fd_sc_hd__inv_1 U161 ( .A(pcgen_icache_va[56]), .Y(n166) );
  sky130_fd_sc_hd__inv_1 U162 ( .A(pcgen_icache_va[39]), .Y(n487) );
  sky130_fd_sc_hd__inv_2 U163 ( .A(n135), .Y(n218) );
  sky130_fd_sc_hd__nor4_1 U164 ( .A(ifu_iu_chgflw_vld), .B(
        icache_pcgen_inst_vld_gate), .C(icache_pcgen_grant_gate), .D(
        btb_xx_chgflw_vld), .Y(n181) );
  sky130_fd_sc_hd__conb_1 U165 ( .LO(n1), .HI(n_Logic1_) );
  sky130_fd_sc_hd__inv_2 U166 ( .A(n137), .Y(n116) );
  sky130_fd_sc_hd__nand2_1 U167 ( .A(n106), .B(n104), .Y(pcgen_pred_flush_vld)
         );
  sky130_fd_sc_hd__nand2_1 U168 ( .A(n108), .B(n28), .Y(n533) );
  sky130_fd_sc_hd__inv_1 U169 ( .A(pcgen_top_buf_chgflw), .Y(n488) );
  sky130_fd_sc_hd__nand4b_1 U170 ( .A_N(iu_ifu_tar_pc_vld_gate), .B(n488), .C(
        n180), .D(n181), .Y(pcgen_icg_en) );
  sky130_fd_sc_hd__nand2_1 U171 ( .A(pred_pcgen_curflw_vld), .B(n488), .Y(n111) );
  sky130_fd_sc_hd__nand2_1 U172 ( .A(btb_xx_chgflw_vld), .B(n488), .Y(n112) );
  sky130_fd_sc_hd__nand2_1 U173 ( .A(n112), .B(n111), .Y(n219) );
  sky130_fd_sc_hd__a222oi_1 U174 ( .A1(pred_pcgen_curflw_pc[0]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[0]), .B2(n68), .C1(pcgen_ifpc_0), .C2(n62), .Y(
        n107) );
  sky130_fd_sc_hd__inv_1 U175 ( .A(n107), .Y(pcgen_btb_ifpc[0]) );
  sky130_fd_sc_hd__nand2_1 U176 ( .A(n31), .B(n108), .Y(n109) );
  sky130_fd_sc_hd__a222oi_1 U177 ( .A1(rtu_ifu_chgflw_pc[0]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[0]), .B2(n26), .C1(
        pred_pcgen_chgflw_pc[0]), .C2(n71), .Y(n110) );
  sky130_fd_sc_hd__inv_1 U178 ( .A(n110), .Y(ifu_iu_chgflw_pc[0]) );
  sky130_fd_sc_hd__nand4_1 U179 ( .A(n29), .B(n112), .C(n52), .D(n124), .Y(
        n223) );
  sky130_fd_sc_hd__inv_1 U180 ( .A(pcgen_ifpc_0), .Y(n123) );
  sky130_fd_sc_hd__mux2i_1 U181 ( .A0(ifu_iu_chgflw_pc[0]), .A1(
        cp0_xx_mrvbr[0]), .S(n94), .Y(n122) );
  sky130_fd_sc_hd__nand2_1 U182 ( .A(n114), .B(n101), .Y(n119) );
  sky130_fd_sc_hd__a22oi_1 U183 ( .A1(pcgen_btb_ifpc[0]), .A2(n18), .B1(
        icache_pcgen_addr[0]), .B2(n84), .Y(n121) );
  sky130_fd_sc_hd__o211ai_1 U184 ( .A1(n39), .A2(n123), .B1(n122), .C1(n121), 
        .Y(N22) );
  sky130_fd_sc_hd__inv_1 U185 ( .A(cp0_xx_mrvbr[0]), .Y(n126) );
  sky130_fd_sc_hd__nand2_1 U186 ( .A(n101), .B(n124), .Y(n485) );
  sky130_fd_sc_hd__nand2_1 U187 ( .A(n485), .B(n101), .Y(n486) );
  sky130_fd_sc_hd__a22oi_1 U188 ( .A1(n92), .A2(pcgen_btb_ifpc[0]), .B1(
        pcgen_pred_ifpc[0]), .B2(n27), .Y(n125) );
  sky130_fd_sc_hd__o21ai_1 U189 ( .A1(n100), .A2(n126), .B1(n125), .Y(n433) );
  sky130_fd_sc_hd__a222oi_1 U190 ( .A1(pred_pcgen_curflw_pc[1]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[1]), .B2(n67), .C1(pcgen_ifpc_1), .C2(n62), .Y(
        n127) );
  sky130_fd_sc_hd__inv_1 U191 ( .A(n127), .Y(pcgen_btb_ifpc[1]) );
  sky130_fd_sc_hd__a222oi_1 U192 ( .A1(rtu_ifu_chgflw_pc[1]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[1]), .B2(n77), .C1(
        pred_pcgen_chgflw_pc[1]), .C2(n74), .Y(n128) );
  sky130_fd_sc_hd__inv_1 U193 ( .A(n128), .Y(ifu_iu_chgflw_pc[1]) );
  sky130_fd_sc_hd__inv_1 U194 ( .A(pcgen_ifpc_1), .Y(n131) );
  sky130_fd_sc_hd__mux2i_1 U195 ( .A0(ifu_iu_chgflw_pc[1]), .A1(
        cp0_xx_mrvbr[1]), .S(n96), .Y(n130) );
  sky130_fd_sc_hd__a22oi_1 U196 ( .A1(pcgen_btb_ifpc[1]), .A2(n18), .B1(
        icache_pcgen_addr[1]), .B2(n84), .Y(n129) );
  sky130_fd_sc_hd__o211ai_1 U197 ( .A1(n39), .A2(n131), .B1(n130), .C1(n129), 
        .Y(N23) );
  sky130_fd_sc_hd__inv_1 U198 ( .A(cp0_xx_mrvbr[1]), .Y(n133) );
  sky130_fd_sc_hd__a22oi_1 U199 ( .A1(n93), .A2(pcgen_btb_ifpc[1]), .B1(
        pcgen_pred_ifpc[1]), .B2(n27), .Y(n132) );
  sky130_fd_sc_hd__o21ai_1 U200 ( .A1(n100), .A2(n133), .B1(n132), .Y(n434) );
  sky130_fd_sc_hd__a222oi_1 U201 ( .A1(pred_pcgen_curflw_pc[2]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[2]), .B2(n67), .C1(pcgen_ifpc_2), .C2(n62), .Y(
        n134) );
  sky130_fd_sc_hd__inv_1 U202 ( .A(n134), .Y(pcgen_btb_ifpc[2]) );
  sky130_fd_sc_hd__inv_1 U203 ( .A(pcgen_ifpc[63]), .Y(n136) );
  sky130_fd_sc_hd__a22o_1 U204 ( .A1(btb_pcgen_tar_pc[39]), .A2(n67), .B1(
        pred_pcgen_curflw_pc[39]), .B2(n69), .X(n135) );
  sky130_fd_sc_hd__o21ai_1 U205 ( .A1(n65), .A2(n136), .B1(n218), .Y(
        pcgen_icache_va[63]) );
  sky130_fd_sc_hd__o21ai_1 U206 ( .A1(n56), .A2(n50), .B1(n97), .Y(n140) );
  sky130_fd_sc_hd__nand2_1 U207 ( .A(n137), .B(icache_pcgen_addr[39]), .Y(n138) );
  sky130_fd_sc_hd__nand2_1 U208 ( .A(n140), .B(n138), .Y(n142) );
  sky130_fd_sc_hd__nand2_1 U209 ( .A(n140), .B(n139), .Y(n141) );
  sky130_fd_sc_hd__nand2_1 U210 ( .A(n142), .B(n141), .Y(n216) );
  sky130_fd_sc_hd__a222oi_1 U211 ( .A1(pcgen_ifpc[63]), .A2(n85), .B1(
        iu_ifu_tar_pc[63]), .B2(n2), .C1(pcgen_ifpc_inc[63]), .C2(n79), .Y(
        n144) );
  sky130_fd_sc_hd__o211ai_1 U212 ( .A1(n30), .A2(n145), .B1(n59), .C1(n144), 
        .Y(N108) );
  sky130_fd_sc_hd__inv_1 U213 ( .A(pcgen_ifpc[62]), .Y(n146) );
  sky130_fd_sc_hd__o21ai_1 U214 ( .A1(n65), .A2(n146), .B1(n218), .Y(
        pcgen_icache_va[62]) );
  sky130_fd_sc_hd__a222oi_1 U215 ( .A1(pcgen_ifpc[62]), .A2(n85), .B1(
        iu_ifu_tar_pc[62]), .B2(n2), .C1(pcgen_ifpc_inc[62]), .C2(n79), .Y(
        n147) );
  sky130_fd_sc_hd__o211ai_1 U216 ( .A1(n30), .A2(n148), .B1(n59), .C1(n147), 
        .Y(N107) );
  sky130_fd_sc_hd__inv_1 U217 ( .A(pcgen_ifpc[61]), .Y(n149) );
  sky130_fd_sc_hd__o21ai_1 U218 ( .A1(n65), .A2(n149), .B1(n218), .Y(
        pcgen_icache_va[61]) );
  sky130_fd_sc_hd__a222oi_1 U219 ( .A1(pcgen_ifpc[61]), .A2(n85), .B1(
        iu_ifu_tar_pc[61]), .B2(n2), .C1(pcgen_ifpc_inc[61]), .C2(n32), .Y(
        n150) );
  sky130_fd_sc_hd__o211ai_1 U220 ( .A1(n30), .A2(n151), .B1(n59), .C1(n150), 
        .Y(N106) );
  sky130_fd_sc_hd__inv_1 U221 ( .A(pcgen_ifpc[60]), .Y(n152) );
  sky130_fd_sc_hd__o21ai_1 U222 ( .A1(n65), .A2(n152), .B1(n218), .Y(
        pcgen_icache_va[60]) );
  sky130_fd_sc_hd__a222oi_1 U223 ( .A1(pcgen_ifpc[60]), .A2(n85), .B1(
        iu_ifu_tar_pc[60]), .B2(n2), .C1(pcgen_ifpc_inc[60]), .C2(n78), .Y(
        n153) );
  sky130_fd_sc_hd__o211ai_1 U224 ( .A1(n30), .A2(n154), .B1(n59), .C1(n153), 
        .Y(N105) );
  sky130_fd_sc_hd__inv_1 U225 ( .A(pcgen_ifpc[59]), .Y(n155) );
  sky130_fd_sc_hd__o21ai_1 U226 ( .A1(n65), .A2(n155), .B1(n218), .Y(
        pcgen_icache_va[59]) );
  sky130_fd_sc_hd__a222oi_1 U227 ( .A1(pcgen_ifpc[59]), .A2(n85), .B1(
        iu_ifu_tar_pc[59]), .B2(n2), .C1(pcgen_ifpc_inc[59]), .C2(n79), .Y(
        n156) );
  sky130_fd_sc_hd__o211ai_1 U228 ( .A1(n30), .A2(n157), .B1(n59), .C1(n156), 
        .Y(N104) );
  sky130_fd_sc_hd__inv_1 U229 ( .A(pcgen_ifpc[58]), .Y(n158) );
  sky130_fd_sc_hd__o21ai_1 U230 ( .A1(n65), .A2(n158), .B1(n218), .Y(
        pcgen_icache_va[58]) );
  sky130_fd_sc_hd__a222oi_1 U231 ( .A1(pcgen_ifpc[58]), .A2(n85), .B1(
        iu_ifu_tar_pc[58]), .B2(n2), .C1(pcgen_ifpc_inc[58]), .C2(n80), .Y(
        n159) );
  sky130_fd_sc_hd__o211ai_1 U232 ( .A1(n30), .A2(n160), .B1(n59), .C1(n159), 
        .Y(N103) );
  sky130_fd_sc_hd__inv_1 U233 ( .A(pcgen_ifpc[57]), .Y(n161) );
  sky130_fd_sc_hd__o21ai_1 U234 ( .A1(n65), .A2(n161), .B1(n218), .Y(
        pcgen_icache_va[57]) );
  sky130_fd_sc_hd__a222oi_1 U235 ( .A1(pcgen_ifpc[57]), .A2(n85), .B1(
        iu_ifu_tar_pc[57]), .B2(n2), .C1(pcgen_ifpc_inc[57]), .C2(n32), .Y(
        n162) );
  sky130_fd_sc_hd__o211ai_1 U236 ( .A1(n30), .A2(n163), .B1(n59), .C1(n162), 
        .Y(N102) );
  sky130_fd_sc_hd__inv_1 U237 ( .A(pcgen_ifpc[56]), .Y(n164) );
  sky130_fd_sc_hd__o21ai_1 U238 ( .A1(n65), .A2(n164), .B1(n218), .Y(
        pcgen_icache_va[56]) );
  sky130_fd_sc_hd__a222oi_1 U239 ( .A1(pcgen_ifpc[56]), .A2(n86), .B1(
        iu_ifu_tar_pc[56]), .B2(n2), .C1(pcgen_ifpc_inc[56]), .C2(n79), .Y(
        n165) );
  sky130_fd_sc_hd__o211ai_1 U240 ( .A1(n30), .A2(n166), .B1(n59), .C1(n165), 
        .Y(N101) );
  sky130_fd_sc_hd__inv_1 U241 ( .A(pcgen_ifpc[55]), .Y(n167) );
  sky130_fd_sc_hd__o21ai_1 U242 ( .A1(n65), .A2(n167), .B1(n218), .Y(
        pcgen_icache_va[55]) );
  sky130_fd_sc_hd__a222oi_1 U243 ( .A1(pcgen_ifpc[55]), .A2(n86), .B1(
        iu_ifu_tar_pc[55]), .B2(n2), .C1(pcgen_ifpc_inc[55]), .C2(n78), .Y(
        n168) );
  sky130_fd_sc_hd__o211ai_1 U244 ( .A1(n30), .A2(n169), .B1(n59), .C1(n168), 
        .Y(N100) );
  sky130_fd_sc_hd__inv_1 U245 ( .A(pcgen_ifpc[54]), .Y(n170) );
  sky130_fd_sc_hd__o21ai_1 U246 ( .A1(n66), .A2(n170), .B1(n218), .Y(
        pcgen_icache_va[54]) );
  sky130_fd_sc_hd__a222oi_1 U247 ( .A1(pcgen_ifpc[54]), .A2(n85), .B1(
        iu_ifu_tar_pc[54]), .B2(n2), .C1(pcgen_ifpc_inc[54]), .C2(n80), .Y(
        n171) );
  sky130_fd_sc_hd__o211ai_1 U248 ( .A1(n30), .A2(n172), .B1(n59), .C1(n171), 
        .Y(N99) );
  sky130_fd_sc_hd__inv_1 U249 ( .A(pcgen_ifpc[53]), .Y(n173) );
  sky130_fd_sc_hd__o21ai_1 U250 ( .A1(n66), .A2(n173), .B1(n218), .Y(
        pcgen_icache_va[53]) );
  sky130_fd_sc_hd__a222oi_1 U251 ( .A1(pcgen_ifpc[53]), .A2(n86), .B1(
        iu_ifu_tar_pc[53]), .B2(n2), .C1(pcgen_ifpc_inc[53]), .C2(n81), .Y(
        n174) );
  sky130_fd_sc_hd__o211ai_1 U252 ( .A1(n30), .A2(n175), .B1(n59), .C1(n174), 
        .Y(N98) );
  sky130_fd_sc_hd__inv_1 U253 ( .A(pcgen_ifpc[52]), .Y(n176) );
  sky130_fd_sc_hd__o21ai_1 U254 ( .A1(n66), .A2(n176), .B1(n218), .Y(
        pcgen_icache_va[52]) );
  sky130_fd_sc_hd__a222oi_1 U255 ( .A1(pcgen_ifpc[52]), .A2(n85), .B1(
        iu_ifu_tar_pc[52]), .B2(n2), .C1(pcgen_ifpc_inc[52]), .C2(n80), .Y(
        n177) );
  sky130_fd_sc_hd__o211ai_1 U256 ( .A1(n30), .A2(n178), .B1(n59), .C1(n177), 
        .Y(N97) );
  sky130_fd_sc_hd__inv_1 U257 ( .A(pcgen_ifpc[51]), .Y(n179) );
  sky130_fd_sc_hd__o21ai_1 U258 ( .A1(n66), .A2(n179), .B1(n218), .Y(
        pcgen_icache_va[51]) );
  sky130_fd_sc_hd__a222oi_1 U259 ( .A1(pcgen_ifpc[51]), .A2(n86), .B1(
        iu_ifu_tar_pc[51]), .B2(n2), .C1(pcgen_ifpc_inc[51]), .C2(n81), .Y(
        n182) );
  sky130_fd_sc_hd__o211ai_1 U260 ( .A1(n30), .A2(n183), .B1(n59), .C1(n182), 
        .Y(N96) );
  sky130_fd_sc_hd__inv_1 U261 ( .A(pcgen_ifpc[50]), .Y(n184) );
  sky130_fd_sc_hd__o21ai_1 U262 ( .A1(n66), .A2(n184), .B1(n218), .Y(
        pcgen_icache_va[50]) );
  sky130_fd_sc_hd__a222oi_1 U263 ( .A1(pcgen_ifpc[50]), .A2(n86), .B1(
        iu_ifu_tar_pc[50]), .B2(n2), .C1(pcgen_ifpc_inc[50]), .C2(n32), .Y(
        n185) );
  sky130_fd_sc_hd__o211ai_1 U264 ( .A1(n30), .A2(n186), .B1(n60), .C1(n185), 
        .Y(N95) );
  sky130_fd_sc_hd__inv_1 U265 ( .A(pcgen_ifpc[49]), .Y(n187) );
  sky130_fd_sc_hd__o21ai_1 U266 ( .A1(n66), .A2(n187), .B1(n218), .Y(
        pcgen_icache_va[49]) );
  sky130_fd_sc_hd__a222oi_1 U267 ( .A1(pcgen_ifpc[49]), .A2(n86), .B1(
        iu_ifu_tar_pc[49]), .B2(n2), .C1(pcgen_ifpc_inc[49]), .C2(n78), .Y(
        n188) );
  sky130_fd_sc_hd__o211ai_1 U268 ( .A1(n30), .A2(n189), .B1(n60), .C1(n188), 
        .Y(N94) );
  sky130_fd_sc_hd__inv_1 U269 ( .A(pcgen_ifpc[48]), .Y(n190) );
  sky130_fd_sc_hd__o21ai_1 U270 ( .A1(n66), .A2(n190), .B1(n218), .Y(
        pcgen_icache_va[48]) );
  sky130_fd_sc_hd__a222oi_1 U271 ( .A1(pcgen_ifpc[48]), .A2(n85), .B1(
        iu_ifu_tar_pc[48]), .B2(n2), .C1(pcgen_ifpc_inc[48]), .C2(n79), .Y(
        n191) );
  sky130_fd_sc_hd__o211ai_1 U272 ( .A1(n30), .A2(n192), .B1(n60), .C1(n191), 
        .Y(N93) );
  sky130_fd_sc_hd__inv_1 U273 ( .A(pcgen_ifpc[47]), .Y(n193) );
  sky130_fd_sc_hd__o21ai_1 U274 ( .A1(n66), .A2(n193), .B1(n218), .Y(
        pcgen_icache_va[47]) );
  sky130_fd_sc_hd__a222oi_1 U275 ( .A1(pcgen_ifpc[47]), .A2(n85), .B1(
        iu_ifu_tar_pc[47]), .B2(n2), .C1(pcgen_ifpc_inc[47]), .C2(n81), .Y(
        n194) );
  sky130_fd_sc_hd__o211ai_1 U276 ( .A1(n30), .A2(n195), .B1(n60), .C1(n194), 
        .Y(N92) );
  sky130_fd_sc_hd__inv_1 U277 ( .A(pcgen_ifpc[46]), .Y(n196) );
  sky130_fd_sc_hd__o21ai_1 U278 ( .A1(n66), .A2(n196), .B1(n218), .Y(
        pcgen_icache_va[46]) );
  sky130_fd_sc_hd__a222oi_1 U279 ( .A1(pcgen_ifpc[46]), .A2(n86), .B1(
        iu_ifu_tar_pc[46]), .B2(n2), .C1(pcgen_ifpc_inc[46]), .C2(n80), .Y(
        n197) );
  sky130_fd_sc_hd__o211ai_1 U280 ( .A1(n30), .A2(n198), .B1(n60), .C1(n197), 
        .Y(N91) );
  sky130_fd_sc_hd__inv_1 U281 ( .A(pcgen_ifpc[45]), .Y(n199) );
  sky130_fd_sc_hd__o21ai_1 U282 ( .A1(n66), .A2(n199), .B1(n218), .Y(
        pcgen_icache_va[45]) );
  sky130_fd_sc_hd__a222oi_1 U283 ( .A1(pcgen_ifpc[45]), .A2(n86), .B1(
        iu_ifu_tar_pc[45]), .B2(n2), .C1(pcgen_ifpc_inc[45]), .C2(n78), .Y(
        n200) );
  sky130_fd_sc_hd__o211ai_1 U284 ( .A1(n30), .A2(n201), .B1(n60), .C1(n200), 
        .Y(N90) );
  sky130_fd_sc_hd__inv_1 U285 ( .A(pcgen_ifpc[44]), .Y(n202) );
  sky130_fd_sc_hd__o21ai_1 U286 ( .A1(n65), .A2(n202), .B1(n218), .Y(
        pcgen_icache_va[44]) );
  sky130_fd_sc_hd__a222oi_1 U287 ( .A1(pcgen_ifpc[44]), .A2(n86), .B1(
        iu_ifu_tar_pc[44]), .B2(n2), .C1(pcgen_ifpc_inc[44]), .C2(n32), .Y(
        n203) );
  sky130_fd_sc_hd__o211ai_1 U288 ( .A1(n30), .A2(n204), .B1(n60), .C1(n203), 
        .Y(N89) );
  sky130_fd_sc_hd__inv_1 U289 ( .A(pcgen_ifpc[43]), .Y(n205) );
  sky130_fd_sc_hd__o21ai_1 U290 ( .A1(n66), .A2(n205), .B1(n218), .Y(
        pcgen_icache_va[43]) );
  sky130_fd_sc_hd__a222oi_1 U291 ( .A1(pcgen_ifpc[43]), .A2(n85), .B1(
        iu_ifu_tar_pc[43]), .B2(n2), .C1(pcgen_ifpc_inc[43]), .C2(n78), .Y(
        n206) );
  sky130_fd_sc_hd__o211ai_1 U292 ( .A1(n30), .A2(n207), .B1(n60), .C1(n206), 
        .Y(N88) );
  sky130_fd_sc_hd__inv_1 U293 ( .A(pcgen_ifpc[42]), .Y(n208) );
  sky130_fd_sc_hd__o21ai_1 U294 ( .A1(n65), .A2(n208), .B1(n218), .Y(
        pcgen_icache_va[42]) );
  sky130_fd_sc_hd__a222oi_1 U295 ( .A1(pcgen_ifpc[42]), .A2(n86), .B1(
        iu_ifu_tar_pc[42]), .B2(n2), .C1(pcgen_ifpc_inc[42]), .C2(n79), .Y(
        n209) );
  sky130_fd_sc_hd__o211ai_1 U296 ( .A1(n30), .A2(n210), .B1(n60), .C1(n209), 
        .Y(N87) );
  sky130_fd_sc_hd__inv_1 U297 ( .A(pcgen_ifpc[41]), .Y(n211) );
  sky130_fd_sc_hd__o21ai_1 U298 ( .A1(n66), .A2(n211), .B1(n218), .Y(
        pcgen_icache_va[41]) );
  sky130_fd_sc_hd__a222oi_1 U299 ( .A1(pcgen_ifpc[41]), .A2(n85), .B1(
        iu_ifu_tar_pc[41]), .B2(n2), .C1(pcgen_ifpc_inc[41]), .C2(n81), .Y(
        n212) );
  sky130_fd_sc_hd__o211ai_1 U300 ( .A1(n30), .A2(n213), .B1(n60), .C1(n212), 
        .Y(N86) );
  sky130_fd_sc_hd__inv_1 U301 ( .A(pcgen_ifpc[40]), .Y(n214) );
  sky130_fd_sc_hd__o21ai_1 U302 ( .A1(n66), .A2(n214), .B1(n218), .Y(
        pcgen_icache_va[40]) );
  sky130_fd_sc_hd__a222oi_1 U303 ( .A1(pcgen_ifpc[40]), .A2(n85), .B1(
        iu_ifu_tar_pc[40]), .B2(n2), .C1(pcgen_ifpc_inc[40]), .C2(n32), .Y(
        n215) );
  sky130_fd_sc_hd__o211ai_1 U304 ( .A1(n30), .A2(n217), .B1(n60), .C1(n215), 
        .Y(N85) );
  sky130_fd_sc_hd__inv_1 U305 ( .A(pcgen_btb_ifpc[39]), .Y(n224) );
  sky130_fd_sc_hd__o21ai_1 U306 ( .A1(n65), .A2(n224), .B1(n218), .Y(
        pcgen_icache_va[39]) );
  sky130_fd_sc_hd__a211o_1 U307 ( .A1(iu_ifu_tar_pc[39]), .A2(n26), .B1(n50), 
        .C1(n56), .X(ifu_iu_chgflw_pc[39]) );
  sky130_fd_sc_hd__nand2_1 U308 ( .A(cp0_xx_mrvbr[39]), .B(n95), .Y(n483) );
  sky130_fd_sc_hd__a221oi_1 U309 ( .A1(icache_pcgen_addr[39]), .A2(n49), .B1(
        ifu_iu_chgflw_pc[39]), .B2(n99), .C1(n220), .Y(n222) );
  sky130_fd_sc_hd__a22oi_1 U310 ( .A1(pcgen_ifpc_inc[39]), .A2(n81), .B1(n18), 
        .B2(pcgen_icache_va[39]), .Y(n221) );
  sky130_fd_sc_hd__o211ai_1 U311 ( .A1(n224), .A2(n39), .B1(n222), .C1(n221), 
        .Y(N61) );
  sky130_fd_sc_hd__a222oi_1 U312 ( .A1(pred_pcgen_curflw_pc[38]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[38]), .B2(n67), .C1(pcgen_btb_ifpc[38]), .C2(n62), 
        .Y(n225) );
  sky130_fd_sc_hd__inv_1 U313 ( .A(n225), .Y(pcgen_icache_va[38]) );
  sky130_fd_sc_hd__a222oi_1 U314 ( .A1(rtu_ifu_chgflw_pc[38]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[38]), .B2(n76), .C1(
        pred_pcgen_chgflw_pc[38]), .C2(n71), .Y(n226) );
  sky130_fd_sc_hd__inv_1 U315 ( .A(n226), .Y(ifu_iu_chgflw_pc[38]) );
  sky130_fd_sc_hd__inv_1 U316 ( .A(cp0_xx_mrvbr[38]), .Y(n482) );
  sky130_fd_sc_hd__mux2i_1 U317 ( .A0(n226), .A1(n482), .S(n96), .Y(n227) );
  sky130_fd_sc_hd__a221o_1 U318 ( .A1(pcgen_ifpc_inc[38]), .A2(n51), .B1(n364), 
        .B2(pcgen_icache_va[38]), .C1(n227), .X(n228) );
  sky130_fd_sc_hd__a221o_1 U319 ( .A1(n87), .A2(pcgen_btb_ifpc[38]), .B1(
        icache_pcgen_addr[38]), .B2(n82), .C1(n228), .X(N60) );
  sky130_fd_sc_hd__a222oi_1 U320 ( .A1(pred_pcgen_curflw_pc[37]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[37]), .B2(n67), .C1(pcgen_btb_ifpc[37]), .C2(n62), 
        .Y(n229) );
  sky130_fd_sc_hd__inv_1 U321 ( .A(n229), .Y(pcgen_icache_va[37]) );
  sky130_fd_sc_hd__a222oi_1 U322 ( .A1(rtu_ifu_chgflw_pc[37]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[37]), .B2(n76), .C1(
        pred_pcgen_chgflw_pc[37]), .C2(n74), .Y(n230) );
  sky130_fd_sc_hd__inv_1 U323 ( .A(n230), .Y(ifu_iu_chgflw_pc[37]) );
  sky130_fd_sc_hd__inv_1 U324 ( .A(cp0_xx_mrvbr[37]), .Y(n478) );
  sky130_fd_sc_hd__mux2i_1 U325 ( .A0(n230), .A1(n478), .S(n96), .Y(n231) );
  sky130_fd_sc_hd__a221o_1 U326 ( .A1(pcgen_ifpc_inc[37]), .A2(n12), .B1(n364), 
        .B2(pcgen_icache_va[37]), .C1(n231), .X(n232) );
  sky130_fd_sc_hd__a221o_1 U327 ( .A1(n86), .A2(pcgen_btb_ifpc[37]), .B1(
        icache_pcgen_addr[37]), .B2(n82), .C1(n232), .X(N59) );
  sky130_fd_sc_hd__a222oi_1 U328 ( .A1(pred_pcgen_curflw_pc[36]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[36]), .B2(n67), .C1(pcgen_btb_ifpc[36]), .C2(n62), 
        .Y(n233) );
  sky130_fd_sc_hd__inv_1 U329 ( .A(n233), .Y(pcgen_icache_va[36]) );
  sky130_fd_sc_hd__a222oi_1 U330 ( .A1(rtu_ifu_chgflw_pc[36]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[36]), .B2(n77), .C1(
        pred_pcgen_chgflw_pc[36]), .C2(n73), .Y(n234) );
  sky130_fd_sc_hd__inv_1 U331 ( .A(n234), .Y(ifu_iu_chgflw_pc[36]) );
  sky130_fd_sc_hd__inv_1 U332 ( .A(cp0_xx_mrvbr[36]), .Y(n476) );
  sky130_fd_sc_hd__mux2i_1 U333 ( .A0(n234), .A1(n476), .S(n96), .Y(n235) );
  sky130_fd_sc_hd__a221o_1 U334 ( .A1(pcgen_ifpc_inc[36]), .A2(n12), .B1(n364), 
        .B2(pcgen_icache_va[36]), .C1(n235), .X(n236) );
  sky130_fd_sc_hd__a221o_1 U335 ( .A1(n86), .A2(pcgen_btb_ifpc[36]), .B1(
        icache_pcgen_addr[36]), .B2(n82), .C1(n236), .X(N58) );
  sky130_fd_sc_hd__a222oi_1 U336 ( .A1(pred_pcgen_curflw_pc[35]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[35]), .B2(n67), .C1(pcgen_btb_ifpc[35]), .C2(n62), 
        .Y(n237) );
  sky130_fd_sc_hd__inv_1 U337 ( .A(n237), .Y(pcgen_icache_va[35]) );
  sky130_fd_sc_hd__a222oi_1 U338 ( .A1(rtu_ifu_chgflw_pc[35]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[35]), .B2(n25), .C1(
        pred_pcgen_chgflw_pc[35]), .C2(n73), .Y(n238) );
  sky130_fd_sc_hd__inv_1 U339 ( .A(n238), .Y(ifu_iu_chgflw_pc[35]) );
  sky130_fd_sc_hd__inv_1 U340 ( .A(cp0_xx_mrvbr[35]), .Y(n474) );
  sky130_fd_sc_hd__mux2i_1 U341 ( .A0(n238), .A1(n474), .S(n96), .Y(n239) );
  sky130_fd_sc_hd__a221o_1 U342 ( .A1(pcgen_ifpc_inc[35]), .A2(n51), .B1(n364), 
        .B2(pcgen_icache_va[35]), .C1(n239), .X(n240) );
  sky130_fd_sc_hd__a221o_1 U343 ( .A1(n85), .A2(pcgen_btb_ifpc[35]), .B1(
        icache_pcgen_addr[35]), .B2(n82), .C1(n240), .X(N57) );
  sky130_fd_sc_hd__a222oi_1 U344 ( .A1(pred_pcgen_curflw_pc[34]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[34]), .B2(n67), .C1(pcgen_btb_ifpc[34]), .C2(n62), 
        .Y(n241) );
  sky130_fd_sc_hd__inv_1 U345 ( .A(n241), .Y(pcgen_icache_va[34]) );
  sky130_fd_sc_hd__a222oi_1 U346 ( .A1(rtu_ifu_chgflw_pc[34]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[34]), .B2(n26), .C1(
        pred_pcgen_chgflw_pc[34]), .C2(n73), .Y(n242) );
  sky130_fd_sc_hd__inv_1 U347 ( .A(n242), .Y(ifu_iu_chgflw_pc[34]) );
  sky130_fd_sc_hd__inv_1 U348 ( .A(cp0_xx_mrvbr[34]), .Y(n432) );
  sky130_fd_sc_hd__mux2i_1 U349 ( .A0(n242), .A1(n432), .S(n96), .Y(n243) );
  sky130_fd_sc_hd__a221o_1 U350 ( .A1(pcgen_ifpc_inc[34]), .A2(n51), .B1(n364), 
        .B2(pcgen_icache_va[34]), .C1(n243), .X(n244) );
  sky130_fd_sc_hd__a221o_1 U351 ( .A1(n86), .A2(pcgen_btb_ifpc[34]), .B1(
        icache_pcgen_addr[34]), .B2(n82), .C1(n244), .X(N56) );
  sky130_fd_sc_hd__a222oi_1 U352 ( .A1(pred_pcgen_curflw_pc[33]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[33]), .B2(n67), .C1(pcgen_btb_ifpc[33]), .C2(n62), 
        .Y(n245) );
  sky130_fd_sc_hd__inv_1 U353 ( .A(n245), .Y(pcgen_icache_va[33]) );
  sky130_fd_sc_hd__a222oi_1 U354 ( .A1(rtu_ifu_chgflw_pc[33]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[33]), .B2(n76), .C1(
        pred_pcgen_chgflw_pc[33]), .C2(n73), .Y(n246) );
  sky130_fd_sc_hd__inv_1 U355 ( .A(n246), .Y(ifu_iu_chgflw_pc[33]) );
  sky130_fd_sc_hd__inv_1 U356 ( .A(cp0_xx_mrvbr[33]), .Y(n430) );
  sky130_fd_sc_hd__mux2i_1 U357 ( .A0(n246), .A1(n430), .S(n96), .Y(n247) );
  sky130_fd_sc_hd__a221o_1 U358 ( .A1(pcgen_ifpc_inc[33]), .A2(n51), .B1(n364), 
        .B2(pcgen_icache_va[33]), .C1(n247), .X(n248) );
  sky130_fd_sc_hd__a221o_1 U359 ( .A1(n87), .A2(pcgen_btb_ifpc[33]), .B1(
        icache_pcgen_addr[33]), .B2(n82), .C1(n248), .X(N55) );
  sky130_fd_sc_hd__a222oi_1 U360 ( .A1(pred_pcgen_curflw_pc[32]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[32]), .B2(n67), .C1(pcgen_btb_ifpc[32]), .C2(n62), 
        .Y(n249) );
  sky130_fd_sc_hd__inv_1 U361 ( .A(n249), .Y(pcgen_icache_va[32]) );
  sky130_fd_sc_hd__a222oi_1 U362 ( .A1(rtu_ifu_chgflw_pc[32]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[32]), .B2(n76), .C1(
        pred_pcgen_chgflw_pc[32]), .C2(n73), .Y(n250) );
  sky130_fd_sc_hd__inv_1 U363 ( .A(n250), .Y(ifu_iu_chgflw_pc[32]) );
  sky130_fd_sc_hd__inv_1 U364 ( .A(cp0_xx_mrvbr[32]), .Y(n428) );
  sky130_fd_sc_hd__mux2i_1 U365 ( .A0(n250), .A1(n428), .S(n96), .Y(n251) );
  sky130_fd_sc_hd__a221o_1 U366 ( .A1(pcgen_ifpc_inc[32]), .A2(n12), .B1(n364), 
        .B2(pcgen_icache_va[32]), .C1(n251), .X(n252) );
  sky130_fd_sc_hd__a221o_1 U367 ( .A1(n86), .A2(pcgen_btb_ifpc[32]), .B1(
        icache_pcgen_addr[32]), .B2(n82), .C1(n252), .X(N54) );
  sky130_fd_sc_hd__a222oi_1 U368 ( .A1(pred_pcgen_curflw_pc[31]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[31]), .B2(n67), .C1(pcgen_btb_ifpc[31]), .C2(n62), 
        .Y(n253) );
  sky130_fd_sc_hd__inv_1 U369 ( .A(n253), .Y(pcgen_icache_va[31]) );
  sky130_fd_sc_hd__a222oi_1 U370 ( .A1(rtu_ifu_chgflw_pc[31]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[31]), .B2(n77), .C1(
        pred_pcgen_chgflw_pc[31]), .C2(n71), .Y(n254) );
  sky130_fd_sc_hd__inv_1 U371 ( .A(n254), .Y(ifu_iu_chgflw_pc[31]) );
  sky130_fd_sc_hd__inv_1 U372 ( .A(cp0_xx_mrvbr[31]), .Y(n426) );
  sky130_fd_sc_hd__mux2i_1 U373 ( .A0(n254), .A1(n426), .S(n96), .Y(n255) );
  sky130_fd_sc_hd__a221o_1 U374 ( .A1(pcgen_ifpc_inc[31]), .A2(n12), .B1(n364), 
        .B2(pcgen_icache_va[31]), .C1(n255), .X(n256) );
  sky130_fd_sc_hd__a221o_1 U375 ( .A1(n86), .A2(pcgen_btb_ifpc[31]), .B1(
        icache_pcgen_addr[31]), .B2(n83), .C1(n256), .X(N53) );
  sky130_fd_sc_hd__a222oi_1 U376 ( .A1(pred_pcgen_curflw_pc[30]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[30]), .B2(n67), .C1(pcgen_btb_ifpc[30]), .C2(n62), 
        .Y(n257) );
  sky130_fd_sc_hd__inv_1 U377 ( .A(n257), .Y(pcgen_icache_va[30]) );
  sky130_fd_sc_hd__a222oi_1 U378 ( .A1(rtu_ifu_chgflw_pc[30]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[30]), .B2(n25), .C1(
        pred_pcgen_chgflw_pc[30]), .C2(n74), .Y(n258) );
  sky130_fd_sc_hd__inv_1 U379 ( .A(n258), .Y(ifu_iu_chgflw_pc[30]) );
  sky130_fd_sc_hd__inv_1 U380 ( .A(cp0_xx_mrvbr[30]), .Y(n424) );
  sky130_fd_sc_hd__mux2i_1 U381 ( .A0(n258), .A1(n424), .S(n96), .Y(n259) );
  sky130_fd_sc_hd__a221o_1 U382 ( .A1(pcgen_ifpc_inc[30]), .A2(n51), .B1(n364), 
        .B2(pcgen_icache_va[30]), .C1(n259), .X(n260) );
  sky130_fd_sc_hd__a221o_1 U383 ( .A1(n86), .A2(pcgen_btb_ifpc[30]), .B1(
        icache_pcgen_addr[30]), .B2(n82), .C1(n260), .X(N52) );
  sky130_fd_sc_hd__a222oi_1 U384 ( .A1(pred_pcgen_curflw_pc[29]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[29]), .B2(n67), .C1(pcgen_btb_ifpc[29]), .C2(n62), 
        .Y(n261) );
  sky130_fd_sc_hd__inv_1 U385 ( .A(n261), .Y(pcgen_icache_va[29]) );
  sky130_fd_sc_hd__a222oi_1 U386 ( .A1(rtu_ifu_chgflw_pc[29]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[29]), .B2(n76), .C1(
        pred_pcgen_chgflw_pc[29]), .C2(n73), .Y(n262) );
  sky130_fd_sc_hd__inv_1 U387 ( .A(n262), .Y(ifu_iu_chgflw_pc[29]) );
  sky130_fd_sc_hd__inv_1 U388 ( .A(cp0_xx_mrvbr[29]), .Y(n422) );
  sky130_fd_sc_hd__mux2i_1 U389 ( .A0(n262), .A1(n422), .S(n96), .Y(n263) );
  sky130_fd_sc_hd__a221o_1 U390 ( .A1(pcgen_ifpc_inc[29]), .A2(n12), .B1(n364), 
        .B2(pcgen_icache_va[29]), .C1(n263), .X(n264) );
  sky130_fd_sc_hd__a221o_1 U391 ( .A1(n85), .A2(pcgen_btb_ifpc[29]), .B1(
        icache_pcgen_addr[29]), .B2(n82), .C1(n264), .X(N51) );
  sky130_fd_sc_hd__a222oi_1 U392 ( .A1(pred_pcgen_curflw_pc[28]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[28]), .B2(n68), .C1(pcgen_btb_ifpc[28]), .C2(n62), 
        .Y(n265) );
  sky130_fd_sc_hd__inv_1 U393 ( .A(n265), .Y(pcgen_icache_va[28]) );
  sky130_fd_sc_hd__a222oi_1 U394 ( .A1(rtu_ifu_chgflw_pc[28]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[28]), .B2(n76), .C1(
        pred_pcgen_chgflw_pc[28]), .C2(n71), .Y(n266) );
  sky130_fd_sc_hd__inv_1 U395 ( .A(n266), .Y(ifu_iu_chgflw_pc[28]) );
  sky130_fd_sc_hd__inv_1 U396 ( .A(cp0_xx_mrvbr[28]), .Y(n420) );
  sky130_fd_sc_hd__mux2i_1 U397 ( .A0(n266), .A1(n420), .S(n96), .Y(n267) );
  sky130_fd_sc_hd__a221o_1 U398 ( .A1(pcgen_ifpc_inc[28]), .A2(n51), .B1(n364), 
        .B2(pcgen_icache_va[28]), .C1(n267), .X(n268) );
  sky130_fd_sc_hd__a221o_1 U399 ( .A1(n86), .A2(pcgen_btb_ifpc[28]), .B1(
        icache_pcgen_addr[28]), .B2(n82), .C1(n268), .X(N50) );
  sky130_fd_sc_hd__a222oi_1 U400 ( .A1(pred_pcgen_curflw_pc[27]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[27]), .B2(n68), .C1(pcgen_btb_ifpc[27]), .C2(n62), 
        .Y(n269) );
  sky130_fd_sc_hd__inv_1 U401 ( .A(n269), .Y(pcgen_icache_va[27]) );
  sky130_fd_sc_hd__a222oi_1 U402 ( .A1(rtu_ifu_chgflw_pc[27]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[27]), .B2(n77), .C1(
        pred_pcgen_chgflw_pc[27]), .C2(n74), .Y(n270) );
  sky130_fd_sc_hd__inv_1 U403 ( .A(n270), .Y(ifu_iu_chgflw_pc[27]) );
  sky130_fd_sc_hd__inv_1 U404 ( .A(cp0_xx_mrvbr[27]), .Y(n418) );
  sky130_fd_sc_hd__mux2i_1 U405 ( .A0(n270), .A1(n418), .S(n96), .Y(n271) );
  sky130_fd_sc_hd__a221o_1 U406 ( .A1(pcgen_ifpc_inc[27]), .A2(n12), .B1(n364), 
        .B2(pcgen_icache_va[27]), .C1(n271), .X(n272) );
  sky130_fd_sc_hd__a221o_1 U407 ( .A1(n87), .A2(pcgen_btb_ifpc[27]), .B1(
        icache_pcgen_addr[27]), .B2(n82), .C1(n272), .X(N49) );
  sky130_fd_sc_hd__a222oi_1 U408 ( .A1(pred_pcgen_curflw_pc[26]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[26]), .B2(n68), .C1(pcgen_btb_ifpc[26]), .C2(n62), 
        .Y(n273) );
  sky130_fd_sc_hd__inv_1 U409 ( .A(n273), .Y(pcgen_icache_va[26]) );
  sky130_fd_sc_hd__a222oi_1 U410 ( .A1(rtu_ifu_chgflw_pc[26]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[26]), .B2(n25), .C1(
        pred_pcgen_chgflw_pc[26]), .C2(n72), .Y(n274) );
  sky130_fd_sc_hd__inv_1 U411 ( .A(n274), .Y(ifu_iu_chgflw_pc[26]) );
  sky130_fd_sc_hd__inv_1 U412 ( .A(cp0_xx_mrvbr[26]), .Y(n416) );
  sky130_fd_sc_hd__mux2i_1 U413 ( .A0(n274), .A1(n416), .S(n95), .Y(n275) );
  sky130_fd_sc_hd__a221o_1 U414 ( .A1(pcgen_ifpc_inc[26]), .A2(n12), .B1(n364), 
        .B2(pcgen_icache_va[26]), .C1(n275), .X(n276) );
  sky130_fd_sc_hd__a221o_1 U415 ( .A1(n86), .A2(pcgen_btb_ifpc[26]), .B1(
        icache_pcgen_addr[26]), .B2(n82), .C1(n276), .X(N48) );
  sky130_fd_sc_hd__a222oi_1 U416 ( .A1(pred_pcgen_curflw_pc[25]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[25]), .B2(n68), .C1(pcgen_btb_ifpc[25]), .C2(n62), 
        .Y(n277) );
  sky130_fd_sc_hd__inv_1 U417 ( .A(n277), .Y(pcgen_icache_va[25]) );
  sky130_fd_sc_hd__a222oi_1 U418 ( .A1(rtu_ifu_chgflw_pc[25]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[25]), .B2(n26), .C1(
        pred_pcgen_chgflw_pc[25]), .C2(n72), .Y(n278) );
  sky130_fd_sc_hd__inv_1 U419 ( .A(n278), .Y(ifu_iu_chgflw_pc[25]) );
  sky130_fd_sc_hd__inv_1 U420 ( .A(cp0_xx_mrvbr[25]), .Y(n414) );
  sky130_fd_sc_hd__mux2i_1 U421 ( .A0(n278), .A1(n414), .S(n95), .Y(n279) );
  sky130_fd_sc_hd__a221o_1 U422 ( .A1(pcgen_ifpc_inc[25]), .A2(n51), .B1(n364), 
        .B2(pcgen_icache_va[25]), .C1(n279), .X(n280) );
  sky130_fd_sc_hd__a221o_1 U423 ( .A1(n86), .A2(pcgen_btb_ifpc[25]), .B1(
        icache_pcgen_addr[25]), .B2(n83), .C1(n280), .X(N47) );
  sky130_fd_sc_hd__a222oi_1 U424 ( .A1(pred_pcgen_curflw_pc[24]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[24]), .B2(n68), .C1(pcgen_btb_ifpc[24]), .C2(n62), 
        .Y(n281) );
  sky130_fd_sc_hd__inv_1 U425 ( .A(n281), .Y(pcgen_icache_va[24]) );
  sky130_fd_sc_hd__a222oi_1 U426 ( .A1(rtu_ifu_chgflw_pc[24]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[24]), .B2(n76), .C1(
        pred_pcgen_chgflw_pc[24]), .C2(n72), .Y(n282) );
  sky130_fd_sc_hd__inv_1 U427 ( .A(n282), .Y(ifu_iu_chgflw_pc[24]) );
  sky130_fd_sc_hd__inv_1 U428 ( .A(cp0_xx_mrvbr[24]), .Y(n412) );
  sky130_fd_sc_hd__mux2i_1 U429 ( .A0(n282), .A1(n412), .S(n95), .Y(n283) );
  sky130_fd_sc_hd__a221o_1 U430 ( .A1(pcgen_ifpc_inc[24]), .A2(n12), .B1(n364), 
        .B2(pcgen_icache_va[24]), .C1(n283), .X(n284) );
  sky130_fd_sc_hd__a221o_1 U431 ( .A1(n85), .A2(pcgen_btb_ifpc[24]), .B1(
        icache_pcgen_addr[24]), .B2(n83), .C1(n284), .X(N46) );
  sky130_fd_sc_hd__a222oi_1 U432 ( .A1(pred_pcgen_curflw_pc[23]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[23]), .B2(n68), .C1(pcgen_btb_ifpc[23]), .C2(n62), 
        .Y(n285) );
  sky130_fd_sc_hd__inv_1 U433 ( .A(n285), .Y(pcgen_icache_va[23]) );
  sky130_fd_sc_hd__a222oi_1 U434 ( .A1(rtu_ifu_chgflw_pc[23]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[23]), .B2(n76), .C1(
        pred_pcgen_chgflw_pc[23]), .C2(n72), .Y(n286) );
  sky130_fd_sc_hd__inv_1 U435 ( .A(n286), .Y(ifu_iu_chgflw_pc[23]) );
  sky130_fd_sc_hd__inv_1 U436 ( .A(cp0_xx_mrvbr[23]), .Y(n410) );
  sky130_fd_sc_hd__mux2i_1 U437 ( .A0(n286), .A1(n410), .S(n95), .Y(n287) );
  sky130_fd_sc_hd__a221o_1 U438 ( .A1(pcgen_ifpc_inc[23]), .A2(n51), .B1(n364), 
        .B2(pcgen_icache_va[23]), .C1(n287), .X(n288) );
  sky130_fd_sc_hd__a221o_1 U439 ( .A1(n86), .A2(pcgen_btb_ifpc[23]), .B1(
        icache_pcgen_addr[23]), .B2(n83), .C1(n288), .X(N45) );
  sky130_fd_sc_hd__a222oi_1 U440 ( .A1(pred_pcgen_curflw_pc[22]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[22]), .B2(n68), .C1(pcgen_btb_ifpc[22]), .C2(n62), 
        .Y(n289) );
  sky130_fd_sc_hd__inv_1 U441 ( .A(n289), .Y(pcgen_icache_va[22]) );
  sky130_fd_sc_hd__a222oi_1 U442 ( .A1(rtu_ifu_chgflw_pc[22]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[22]), .B2(n77), .C1(
        pred_pcgen_chgflw_pc[22]), .C2(n72), .Y(n290) );
  sky130_fd_sc_hd__inv_1 U443 ( .A(n290), .Y(ifu_iu_chgflw_pc[22]) );
  sky130_fd_sc_hd__inv_1 U444 ( .A(cp0_xx_mrvbr[22]), .Y(n408) );
  sky130_fd_sc_hd__mux2i_1 U445 ( .A0(n290), .A1(n408), .S(n95), .Y(n291) );
  sky130_fd_sc_hd__a221o_1 U446 ( .A1(pcgen_ifpc_inc[22]), .A2(n51), .B1(n18), 
        .B2(pcgen_icache_va[22]), .C1(n291), .X(n292) );
  sky130_fd_sc_hd__a221o_1 U447 ( .A1(n87), .A2(pcgen_btb_ifpc[22]), .B1(
        icache_pcgen_addr[22]), .B2(n83), .C1(n292), .X(N44) );
  sky130_fd_sc_hd__a222oi_1 U448 ( .A1(pred_pcgen_curflw_pc[21]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[21]), .B2(n68), .C1(pcgen_btb_ifpc[21]), .C2(n62), 
        .Y(n293) );
  sky130_fd_sc_hd__inv_1 U449 ( .A(n293), .Y(pcgen_icache_va[21]) );
  sky130_fd_sc_hd__a222oi_1 U450 ( .A1(rtu_ifu_chgflw_pc[21]), .A2(
        ifu_iu_chgflw_vld), .B1(iu_ifu_tar_pc[21]), .B2(n25), .C1(
        pred_pcgen_chgflw_pc[21]), .C2(n72), .Y(n294) );
  sky130_fd_sc_hd__inv_1 U451 ( .A(n294), .Y(ifu_iu_chgflw_pc[21]) );
  sky130_fd_sc_hd__inv_1 U452 ( .A(cp0_xx_mrvbr[21]), .Y(n406) );
  sky130_fd_sc_hd__mux2i_1 U453 ( .A0(n294), .A1(n406), .S(n95), .Y(n295) );
  sky130_fd_sc_hd__a221o_1 U454 ( .A1(pcgen_ifpc_inc[21]), .A2(n51), .B1(n18), 
        .B2(pcgen_icache_va[21]), .C1(n295), .X(n296) );
  sky130_fd_sc_hd__a221o_1 U455 ( .A1(n86), .A2(pcgen_btb_ifpc[21]), .B1(
        icache_pcgen_addr[21]), .B2(n83), .C1(n296), .X(N43) );
  sky130_fd_sc_hd__a222oi_1 U456 ( .A1(pred_pcgen_curflw_pc[20]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[20]), .B2(n68), .C1(pcgen_btb_ifpc[20]), .C2(n62), 
        .Y(n297) );
  sky130_fd_sc_hd__inv_1 U457 ( .A(n297), .Y(pcgen_icache_va[20]) );
  sky130_fd_sc_hd__a222oi_1 U458 ( .A1(rtu_ifu_chgflw_pc[20]), .A2(n57), .B1(
        iu_ifu_tar_pc[20]), .B2(n76), .C1(pred_pcgen_chgflw_pc[20]), .C2(n73), 
        .Y(n298) );
  sky130_fd_sc_hd__inv_1 U459 ( .A(n298), .Y(ifu_iu_chgflw_pc[20]) );
  sky130_fd_sc_hd__inv_1 U460 ( .A(cp0_xx_mrvbr[20]), .Y(n404) );
  sky130_fd_sc_hd__mux2i_1 U461 ( .A0(n298), .A1(n404), .S(n95), .Y(n299) );
  sky130_fd_sc_hd__a221o_1 U462 ( .A1(pcgen_ifpc_inc[20]), .A2(n51), .B1(n18), 
        .B2(pcgen_icache_va[20]), .C1(n299), .X(n300) );
  sky130_fd_sc_hd__a221o_1 U463 ( .A1(n86), .A2(pcgen_btb_ifpc[20]), .B1(
        icache_pcgen_addr[20]), .B2(n83), .C1(n300), .X(N42) );
  sky130_fd_sc_hd__a222oi_1 U464 ( .A1(pred_pcgen_curflw_pc[19]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[19]), .B2(n68), .C1(pcgen_btb_ifpc[19]), .C2(n62), 
        .Y(n301) );
  sky130_fd_sc_hd__inv_1 U465 ( .A(n301), .Y(pcgen_icache_va[19]) );
  sky130_fd_sc_hd__a222oi_1 U466 ( .A1(rtu_ifu_chgflw_pc[19]), .A2(n57), .B1(
        iu_ifu_tar_pc[19]), .B2(n76), .C1(pred_pcgen_chgflw_pc[19]), .C2(n73), 
        .Y(n302) );
  sky130_fd_sc_hd__inv_1 U467 ( .A(n302), .Y(ifu_iu_chgflw_pc[19]) );
  sky130_fd_sc_hd__inv_1 U468 ( .A(cp0_xx_mrvbr[19]), .Y(n402) );
  sky130_fd_sc_hd__mux2i_1 U469 ( .A0(n302), .A1(n402), .S(n95), .Y(n303) );
  sky130_fd_sc_hd__a221o_1 U470 ( .A1(pcgen_ifpc_inc[19]), .A2(n12), .B1(n18), 
        .B2(pcgen_icache_va[19]), .C1(n303), .X(n304) );
  sky130_fd_sc_hd__a221o_1 U471 ( .A1(n85), .A2(pcgen_btb_ifpc[19]), .B1(
        icache_pcgen_addr[19]), .B2(n83), .C1(n304), .X(N41) );
  sky130_fd_sc_hd__a222oi_1 U472 ( .A1(pred_pcgen_curflw_pc[18]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[18]), .B2(n68), .C1(pcgen_btb_ifpc[18]), .C2(n62), 
        .Y(n305) );
  sky130_fd_sc_hd__inv_1 U473 ( .A(n305), .Y(pcgen_icache_va[18]) );
  sky130_fd_sc_hd__a222oi_1 U474 ( .A1(rtu_ifu_chgflw_pc[18]), .A2(n57), .B1(
        iu_ifu_tar_pc[18]), .B2(n77), .C1(pred_pcgen_chgflw_pc[18]), .C2(n73), 
        .Y(n306) );
  sky130_fd_sc_hd__inv_1 U475 ( .A(n306), .Y(ifu_iu_chgflw_pc[18]) );
  sky130_fd_sc_hd__inv_1 U476 ( .A(cp0_xx_mrvbr[18]), .Y(n400) );
  sky130_fd_sc_hd__mux2i_1 U477 ( .A0(n306), .A1(n400), .S(n95), .Y(n307) );
  sky130_fd_sc_hd__a221o_1 U478 ( .A1(pcgen_ifpc_inc[18]), .A2(n12), .B1(n18), 
        .B2(pcgen_icache_va[18]), .C1(n307), .X(n308) );
  sky130_fd_sc_hd__a221o_1 U479 ( .A1(n86), .A2(pcgen_btb_ifpc[18]), .B1(
        icache_pcgen_addr[18]), .B2(n83), .C1(n308), .X(N40) );
  sky130_fd_sc_hd__a222oi_1 U480 ( .A1(pred_pcgen_curflw_pc[17]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[17]), .B2(n68), .C1(pcgen_btb_ifpc[17]), .C2(n62), 
        .Y(n309) );
  sky130_fd_sc_hd__inv_1 U481 ( .A(n309), .Y(pcgen_icache_va[17]) );
  sky130_fd_sc_hd__a222oi_1 U482 ( .A1(rtu_ifu_chgflw_pc[17]), .A2(n57), .B1(
        iu_ifu_tar_pc[17]), .B2(n25), .C1(pred_pcgen_chgflw_pc[17]), .C2(n73), 
        .Y(n310) );
  sky130_fd_sc_hd__inv_1 U483 ( .A(n310), .Y(ifu_iu_chgflw_pc[17]) );
  sky130_fd_sc_hd__inv_1 U484 ( .A(cp0_xx_mrvbr[17]), .Y(n398) );
  sky130_fd_sc_hd__mux2i_1 U485 ( .A0(n310), .A1(n398), .S(n95), .Y(n311) );
  sky130_fd_sc_hd__a221o_1 U486 ( .A1(pcgen_ifpc_inc[17]), .A2(n51), .B1(n18), 
        .B2(pcgen_icache_va[17]), .C1(n311), .X(n312) );
  sky130_fd_sc_hd__a221o_1 U487 ( .A1(n87), .A2(pcgen_btb_ifpc[17]), .B1(
        icache_pcgen_addr[17]), .B2(n83), .C1(n312), .X(N39) );
  sky130_fd_sc_hd__a222oi_1 U488 ( .A1(pred_pcgen_curflw_pc[16]), .A2(n70), 
        .B1(btb_pcgen_tar_pc[16]), .B2(n68), .C1(pcgen_btb_ifpc[16]), .C2(n62), 
        .Y(n313) );
  sky130_fd_sc_hd__inv_1 U489 ( .A(n313), .Y(pcgen_icache_va[16]) );
  sky130_fd_sc_hd__a222oi_1 U490 ( .A1(rtu_ifu_chgflw_pc[16]), .A2(n57), .B1(
        iu_ifu_tar_pc[16]), .B2(n26), .C1(pred_pcgen_chgflw_pc[16]), .C2(n73), 
        .Y(n314) );
  sky130_fd_sc_hd__inv_1 U491 ( .A(n314), .Y(ifu_iu_chgflw_pc[16]) );
  sky130_fd_sc_hd__inv_1 U492 ( .A(cp0_xx_mrvbr[16]), .Y(n396) );
  sky130_fd_sc_hd__mux2i_1 U493 ( .A0(n314), .A1(n396), .S(n95), .Y(n315) );
  sky130_fd_sc_hd__a221o_1 U494 ( .A1(pcgen_ifpc_inc[16]), .A2(n12), .B1(n18), 
        .B2(pcgen_icache_va[16]), .C1(n315), .X(n316) );
  sky130_fd_sc_hd__a221o_1 U495 ( .A1(n86), .A2(pcgen_btb_ifpc[16]), .B1(
        icache_pcgen_addr[16]), .B2(n83), .C1(n316), .X(N38) );
  sky130_fd_sc_hd__a222oi_1 U496 ( .A1(pred_pcgen_curflw_pc[15]), .A2(n70), 
        .B1(btb_pcgen_tar_pc[15]), .B2(n53), .C1(pcgen_icache_seq_tag[9]), 
        .C2(n63), .Y(n317) );
  sky130_fd_sc_hd__inv_1 U497 ( .A(n317), .Y(pcgen_btb_ifpc[15]) );
  sky130_fd_sc_hd__a222oi_1 U498 ( .A1(rtu_ifu_chgflw_pc[15]), .A2(n57), .B1(
        iu_ifu_tar_pc[15]), .B2(n75), .C1(pred_pcgen_chgflw_pc[15]), .C2(n73), 
        .Y(n318) );
  sky130_fd_sc_hd__inv_1 U499 ( .A(n318), .Y(ifu_iu_chgflw_pc[15]) );
  sky130_fd_sc_hd__inv_1 U500 ( .A(cp0_xx_mrvbr[15]), .Y(n394) );
  sky130_fd_sc_hd__mux2i_1 U501 ( .A0(n318), .A1(n394), .S(n95), .Y(n319) );
  sky130_fd_sc_hd__a221o_1 U502 ( .A1(pcgen_ifpc_inc[15]), .A2(n51), .B1(n18), 
        .B2(pcgen_btb_ifpc[15]), .C1(n319), .X(n320) );
  sky130_fd_sc_hd__a221o_1 U503 ( .A1(n85), .A2(pcgen_icache_seq_tag[9]), .B1(
        icache_pcgen_addr[15]), .B2(n83), .C1(n320), .X(N37) );
  sky130_fd_sc_hd__a222oi_1 U504 ( .A1(pred_pcgen_curflw_pc[14]), .A2(n70), 
        .B1(btb_pcgen_tar_pc[14]), .B2(n53), .C1(pcgen_icache_seq_tag[8]), 
        .C2(n63), .Y(n321) );
  sky130_fd_sc_hd__inv_1 U505 ( .A(n321), .Y(pcgen_btb_ifpc[14]) );
  sky130_fd_sc_hd__a222oi_1 U506 ( .A1(rtu_ifu_chgflw_pc[14]), .A2(n57), .B1(
        iu_ifu_tar_pc[14]), .B2(n75), .C1(pred_pcgen_chgflw_pc[14]), .C2(n71), 
        .Y(n322) );
  sky130_fd_sc_hd__inv_1 U507 ( .A(n322), .Y(ifu_iu_chgflw_pc[14]) );
  sky130_fd_sc_hd__inv_1 U508 ( .A(cp0_xx_mrvbr[14]), .Y(n392) );
  sky130_fd_sc_hd__mux2i_1 U509 ( .A0(n322), .A1(n392), .S(n94), .Y(n323) );
  sky130_fd_sc_hd__a221o_1 U510 ( .A1(pcgen_ifpc_inc[14]), .A2(n12), .B1(n18), 
        .B2(pcgen_btb_ifpc[14]), .C1(n323), .X(n324) );
  sky130_fd_sc_hd__a221o_1 U511 ( .A1(n86), .A2(pcgen_icache_seq_tag[8]), .B1(
        icache_pcgen_addr[14]), .B2(n83), .C1(n324), .X(N36) );
  sky130_fd_sc_hd__a222oi_1 U512 ( .A1(pred_pcgen_curflw_pc[13]), .A2(n70), 
        .B1(btb_pcgen_tar_pc[13]), .B2(n53), .C1(pcgen_icache_seq_tag[7]), 
        .C2(n63), .Y(n325) );
  sky130_fd_sc_hd__inv_1 U513 ( .A(n325), .Y(pcgen_btb_ifpc[13]) );
  sky130_fd_sc_hd__a222oi_1 U514 ( .A1(rtu_ifu_chgflw_pc[13]), .A2(n57), .B1(
        iu_ifu_tar_pc[13]), .B2(n75), .C1(pred_pcgen_chgflw_pc[13]), .C2(n74), 
        .Y(n326) );
  sky130_fd_sc_hd__inv_1 U515 ( .A(n326), .Y(ifu_iu_chgflw_pc[13]) );
  sky130_fd_sc_hd__inv_1 U516 ( .A(cp0_xx_mrvbr[13]), .Y(n390) );
  sky130_fd_sc_hd__a221o_1 U517 ( .A1(n86), .A2(pcgen_icache_seq_tag[7]), .B1(
        icache_pcgen_addr[13]), .B2(n84), .C1(n327), .X(N35) );
  sky130_fd_sc_hd__a222oi_1 U518 ( .A1(pred_pcgen_curflw_pc[12]), .A2(n70), 
        .B1(btb_pcgen_tar_pc[12]), .B2(n53), .C1(pcgen_icache_seq_tag[6]), 
        .C2(n63), .Y(n328) );
  sky130_fd_sc_hd__inv_1 U519 ( .A(n328), .Y(pcgen_btb_ifpc[12]) );
  sky130_fd_sc_hd__a222oi_1 U520 ( .A1(rtu_ifu_chgflw_pc[12]), .A2(n57), .B1(
        iu_ifu_tar_pc[12]), .B2(n77), .C1(pred_pcgen_chgflw_pc[12]), .C2(n71), 
        .Y(n329) );
  sky130_fd_sc_hd__inv_1 U521 ( .A(n329), .Y(ifu_iu_chgflw_pc[12]) );
  sky130_fd_sc_hd__inv_1 U522 ( .A(cp0_xx_mrvbr[12]), .Y(n388) );
  sky130_fd_sc_hd__mux2i_1 U523 ( .A0(n329), .A1(n388), .S(n94), .Y(n330) );
  sky130_fd_sc_hd__a222oi_1 U524 ( .A1(pred_pcgen_curflw_pc[11]), .A2(n70), 
        .B1(btb_pcgen_tar_pc[11]), .B2(n53), .C1(pcgen_icache_seq_tag[5]), 
        .C2(n63), .Y(n331) );
  sky130_fd_sc_hd__inv_1 U525 ( .A(n331), .Y(pcgen_btb_ifpc[11]) );
  sky130_fd_sc_hd__a222oi_1 U526 ( .A1(rtu_ifu_chgflw_pc[11]), .A2(n57), .B1(
        iu_ifu_tar_pc[11]), .B2(n75), .C1(pred_pcgen_chgflw_pc[11]), .C2(n73), 
        .Y(n332) );
  sky130_fd_sc_hd__inv_1 U527 ( .A(n332), .Y(ifu_iu_chgflw_pc[11]) );
  sky130_fd_sc_hd__inv_1 U528 ( .A(cp0_xx_mrvbr[11]), .Y(n386) );
  sky130_fd_sc_hd__mux2i_1 U529 ( .A0(n332), .A1(n386), .S(n95), .Y(n333) );
  sky130_fd_sc_hd__a222oi_1 U530 ( .A1(pred_pcgen_curflw_pc[10]), .A2(n70), 
        .B1(btb_pcgen_tar_pc[10]), .B2(n53), .C1(pcgen_icache_seq_tag[4]), 
        .C2(n63), .Y(n334) );
  sky130_fd_sc_hd__inv_1 U531 ( .A(n334), .Y(pcgen_btb_ifpc[10]) );
  sky130_fd_sc_hd__a222oi_1 U532 ( .A1(rtu_ifu_chgflw_pc[10]), .A2(n57), .B1(
        iu_ifu_tar_pc[10]), .B2(n25), .C1(pred_pcgen_chgflw_pc[10]), .C2(n74), 
        .Y(n335) );
  sky130_fd_sc_hd__inv_1 U533 ( .A(n335), .Y(ifu_iu_chgflw_pc[10]) );
  sky130_fd_sc_hd__inv_1 U534 ( .A(cp0_xx_mrvbr[10]), .Y(n384) );
  sky130_fd_sc_hd__mux2i_1 U535 ( .A0(n335), .A1(n384), .S(n94), .Y(n336) );
  sky130_fd_sc_hd__a222oi_1 U536 ( .A1(pred_pcgen_curflw_pc[9]), .A2(n70), 
        .B1(btb_pcgen_tar_pc[9]), .B2(n53), .C1(pcgen_icache_seq_tag[3]), .C2(
        n63), .Y(n337) );
  sky130_fd_sc_hd__inv_1 U537 ( .A(n337), .Y(pcgen_btb_ifpc[9]) );
  sky130_fd_sc_hd__a222oi_1 U538 ( .A1(rtu_ifu_chgflw_pc[9]), .A2(n57), .B1(
        iu_ifu_tar_pc[9]), .B2(n77), .C1(pred_pcgen_chgflw_pc[9]), .C2(n71), 
        .Y(n338) );
  sky130_fd_sc_hd__inv_1 U539 ( .A(n338), .Y(ifu_iu_chgflw_pc[9]) );
  sky130_fd_sc_hd__inv_1 U540 ( .A(cp0_xx_mrvbr[9]), .Y(n382) );
  sky130_fd_sc_hd__mux2i_1 U541 ( .A0(n338), .A1(n382), .S(n94), .Y(n339) );
  sky130_fd_sc_hd__a222oi_1 U542 ( .A1(pred_pcgen_curflw_pc[8]), .A2(n70), 
        .B1(btb_pcgen_tar_pc[8]), .B2(n53), .C1(pcgen_icache_seq_tag[2]), .C2(
        n63), .Y(n340) );
  sky130_fd_sc_hd__inv_1 U543 ( .A(n340), .Y(pcgen_btb_ifpc[8]) );
  sky130_fd_sc_hd__a222oi_1 U544 ( .A1(rtu_ifu_chgflw_pc[8]), .A2(n57), .B1(
        iu_ifu_tar_pc[8]), .B2(n26), .C1(pred_pcgen_chgflw_pc[8]), .C2(n73), 
        .Y(n341) );
  sky130_fd_sc_hd__inv_1 U545 ( .A(n341), .Y(ifu_iu_chgflw_pc[8]) );
  sky130_fd_sc_hd__inv_1 U546 ( .A(cp0_xx_mrvbr[8]), .Y(n380) );
  sky130_fd_sc_hd__mux2i_1 U547 ( .A0(n341), .A1(n380), .S(n94), .Y(n342) );
  sky130_fd_sc_hd__a222oi_1 U548 ( .A1(pred_pcgen_curflw_pc[7]), .A2(n70), 
        .B1(btb_pcgen_tar_pc[7]), .B2(n53), .C1(pcgen_icache_seq_tag[1]), .C2(
        n63), .Y(n343) );
  sky130_fd_sc_hd__inv_1 U549 ( .A(n343), .Y(pcgen_btb_ifpc[7]) );
  sky130_fd_sc_hd__a222oi_1 U550 ( .A1(rtu_ifu_chgflw_pc[7]), .A2(n57), .B1(
        iu_ifu_tar_pc[7]), .B2(n75), .C1(pred_pcgen_chgflw_pc[7]), .C2(n73), 
        .Y(n344) );
  sky130_fd_sc_hd__inv_1 U551 ( .A(n344), .Y(ifu_iu_chgflw_pc[7]) );
  sky130_fd_sc_hd__inv_1 U552 ( .A(cp0_xx_mrvbr[7]), .Y(n378) );
  sky130_fd_sc_hd__mux2i_1 U553 ( .A0(n344), .A1(n378), .S(n94), .Y(n345) );
  sky130_fd_sc_hd__a221o_1 U554 ( .A1(pcgen_ifpc_inc[7]), .A2(n51), .B1(n364), 
        .B2(pcgen_btb_ifpc[7]), .C1(n345), .X(n346) );
  sky130_fd_sc_hd__a221o_1 U555 ( .A1(n87), .A2(pcgen_icache_seq_tag[1]), .B1(
        icache_pcgen_addr[7]), .B2(n84), .C1(n346), .X(N29) );
  sky130_fd_sc_hd__a222oi_1 U556 ( .A1(pred_pcgen_curflw_pc[6]), .A2(n70), 
        .B1(btb_pcgen_tar_pc[6]), .B2(n53), .C1(pcgen_icache_seq_tag[0]), .C2(
        n63), .Y(n347) );
  sky130_fd_sc_hd__inv_1 U557 ( .A(n347), .Y(pcgen_btb_ifpc[6]) );
  sky130_fd_sc_hd__a222oi_1 U558 ( .A1(rtu_ifu_chgflw_pc[6]), .A2(n57), .B1(
        iu_ifu_tar_pc[6]), .B2(n25), .C1(pred_pcgen_chgflw_pc[6]), .C2(n74), 
        .Y(n348) );
  sky130_fd_sc_hd__inv_1 U559 ( .A(n348), .Y(ifu_iu_chgflw_pc[6]) );
  sky130_fd_sc_hd__inv_1 U560 ( .A(cp0_xx_mrvbr[6]), .Y(n376) );
  sky130_fd_sc_hd__mux2i_1 U561 ( .A0(n348), .A1(n376), .S(n94), .Y(n349) );
  sky130_fd_sc_hd__a222oi_1 U562 ( .A1(pred_pcgen_curflw_pc[5]), .A2(n70), 
        .B1(btb_pcgen_tar_pc[5]), .B2(n53), .C1(pcgen_ifpc_5), .C2(n63), .Y(
        n350) );
  sky130_fd_sc_hd__inv_1 U563 ( .A(n350), .Y(pcgen_btb_ifpc[5]) );
  sky130_fd_sc_hd__a222oi_1 U564 ( .A1(rtu_ifu_chgflw_pc[5]), .A2(n57), .B1(
        iu_ifu_tar_pc[5]), .B2(n75), .C1(pred_pcgen_chgflw_pc[5]), .C2(n73), 
        .Y(n351) );
  sky130_fd_sc_hd__inv_1 U565 ( .A(n351), .Y(ifu_iu_chgflw_pc[5]) );
  sky130_fd_sc_hd__inv_1 U566 ( .A(cp0_xx_mrvbr[5]), .Y(n374) );
  sky130_fd_sc_hd__mux2i_1 U567 ( .A0(n351), .A1(n374), .S(n94), .Y(n352) );
  sky130_fd_sc_hd__a222oi_1 U568 ( .A1(pred_pcgen_curflw_pc[4]), .A2(n70), 
        .B1(btb_pcgen_tar_pc[4]), .B2(n68), .C1(pcgen_ifpc_4), .C2(n63), .Y(
        n353) );
  sky130_fd_sc_hd__inv_1 U569 ( .A(n353), .Y(pcgen_btb_ifpc[4]) );
  sky130_fd_sc_hd__a222oi_1 U570 ( .A1(rtu_ifu_chgflw_pc[4]), .A2(n57), .B1(
        iu_ifu_tar_pc[4]), .B2(n75), .C1(pred_pcgen_chgflw_pc[4]), .C2(n73), 
        .Y(n354) );
  sky130_fd_sc_hd__inv_1 U571 ( .A(n354), .Y(ifu_iu_chgflw_pc[4]) );
  sky130_fd_sc_hd__inv_1 U572 ( .A(cp0_xx_mrvbr[4]), .Y(n372) );
  sky130_fd_sc_hd__mux2i_1 U573 ( .A0(n354), .A1(n372), .S(n94), .Y(n355) );
  sky130_fd_sc_hd__a221o_1 U574 ( .A1(pcgen_ifpc_inc[4]), .A2(n12), .B1(n364), 
        .B2(pcgen_btb_ifpc[4]), .C1(n355), .X(n356) );
  sky130_fd_sc_hd__a221o_1 U575 ( .A1(n87), .A2(pcgen_ifpc_4), .B1(
        icache_pcgen_addr[4]), .B2(n84), .C1(n356), .X(N26) );
  sky130_fd_sc_hd__a222oi_1 U576 ( .A1(pred_pcgen_curflw_pc[3]), .A2(n69), 
        .B1(btb_pcgen_tar_pc[3]), .B2(n67), .C1(pcgen_ifpc_3), .C2(n63), .Y(
        n358) );
  sky130_fd_sc_hd__inv_1 U577 ( .A(n358), .Y(pcgen_btb_ifpc[3]) );
  sky130_fd_sc_hd__a222oi_1 U578 ( .A1(rtu_ifu_chgflw_pc[3]), .A2(n57), .B1(
        iu_ifu_tar_pc[3]), .B2(n75), .C1(pred_pcgen_chgflw_pc[3]), .C2(n73), 
        .Y(n359) );
  sky130_fd_sc_hd__inv_1 U579 ( .A(n359), .Y(ifu_iu_chgflw_pc[3]) );
  sky130_fd_sc_hd__inv_1 U580 ( .A(cp0_xx_mrvbr[3]), .Y(n370) );
  sky130_fd_sc_hd__mux2i_1 U581 ( .A0(n359), .A1(n370), .S(n94), .Y(n360) );
  sky130_fd_sc_hd__a222oi_1 U582 ( .A1(rtu_ifu_chgflw_pc[2]), .A2(n57), .B1(
        iu_ifu_tar_pc[2]), .B2(n26), .C1(pred_pcgen_chgflw_pc[2]), .C2(n73), 
        .Y(n362) );
  sky130_fd_sc_hd__inv_1 U583 ( .A(n362), .Y(ifu_iu_chgflw_pc[2]) );
  sky130_fd_sc_hd__inv_1 U584 ( .A(cp0_xx_mrvbr[2]), .Y(n368) );
  sky130_fd_sc_hd__mux2i_1 U585 ( .A0(n362), .A1(n368), .S(n94), .Y(n363) );
  sky130_fd_sc_hd__a221o_1 U586 ( .A1(pcgen_ifpc_inc[2]), .A2(n12), .B1(n18), 
        .B2(pcgen_btb_ifpc[2]), .C1(n363), .X(n365) );
  sky130_fd_sc_hd__a221o_1 U587 ( .A1(n87), .A2(pcgen_ifpc_2), .B1(
        icache_pcgen_addr[2]), .B2(n82), .C1(n365), .X(N24) );
  sky130_fd_sc_hd__a22oi_1 U588 ( .A1(n11), .A2(pcgen_btb_ifpc[2]), .B1(
        pcgen_pred_ifpc[2]), .B2(n90), .Y(n367) );
  sky130_fd_sc_hd__o21ai_1 U589 ( .A1(n100), .A2(n368), .B1(n367), .Y(n435) );
  sky130_fd_sc_hd__a22oi_1 U590 ( .A1(n10), .A2(pcgen_btb_ifpc[3]), .B1(
        pcgen_pred_ifpc[3]), .B2(n89), .Y(n369) );
  sky130_fd_sc_hd__o21ai_1 U591 ( .A1(n100), .A2(n370), .B1(n369), .Y(n436) );
  sky130_fd_sc_hd__a22oi_1 U592 ( .A1(n92), .A2(pcgen_btb_ifpc[4]), .B1(
        pcgen_pred_ifpc[4]), .B2(n27), .Y(n371) );
  sky130_fd_sc_hd__o21ai_1 U593 ( .A1(n100), .A2(n372), .B1(n371), .Y(n437) );
  sky130_fd_sc_hd__a22oi_1 U594 ( .A1(n93), .A2(pcgen_btb_ifpc[5]), .B1(
        pcgen_pred_ifpc[5]), .B2(n27), .Y(n373) );
  sky130_fd_sc_hd__o21ai_1 U595 ( .A1(n100), .A2(n374), .B1(n373), .Y(n438) );
  sky130_fd_sc_hd__a22oi_1 U596 ( .A1(n11), .A2(pcgen_btb_ifpc[6]), .B1(
        pcgen_pred_ifpc[6]), .B2(n27), .Y(n375) );
  sky130_fd_sc_hd__o21ai_1 U597 ( .A1(n100), .A2(n376), .B1(n375), .Y(n439) );
  sky130_fd_sc_hd__a22oi_1 U598 ( .A1(n10), .A2(pcgen_btb_ifpc[7]), .B1(
        pcgen_pred_ifpc[7]), .B2(n27), .Y(n377) );
  sky130_fd_sc_hd__o21ai_1 U599 ( .A1(n100), .A2(n378), .B1(n377), .Y(n440) );
  sky130_fd_sc_hd__a22oi_1 U600 ( .A1(n10), .A2(pcgen_btb_ifpc[8]), .B1(
        pcgen_pred_ifpc[8]), .B2(n89), .Y(n379) );
  sky130_fd_sc_hd__o21ai_1 U601 ( .A1(n99), .A2(n380), .B1(n379), .Y(n441) );
  sky130_fd_sc_hd__a22oi_1 U602 ( .A1(n92), .A2(pcgen_btb_ifpc[9]), .B1(
        pcgen_pred_ifpc[9]), .B2(n27), .Y(n381) );
  sky130_fd_sc_hd__o21ai_1 U603 ( .A1(n99), .A2(n382), .B1(n381), .Y(n442) );
  sky130_fd_sc_hd__a22oi_1 U604 ( .A1(n93), .A2(pcgen_btb_ifpc[10]), .B1(
        pcgen_pred_ifpc[10]), .B2(n27), .Y(n383) );
  sky130_fd_sc_hd__o21ai_1 U605 ( .A1(n99), .A2(n384), .B1(n383), .Y(n443) );
  sky130_fd_sc_hd__a22oi_1 U606 ( .A1(n11), .A2(pcgen_btb_ifpc[11]), .B1(
        pcgen_pred_ifpc[11]), .B2(n90), .Y(n385) );
  sky130_fd_sc_hd__o21ai_1 U607 ( .A1(n99), .A2(n386), .B1(n385), .Y(n444) );
  sky130_fd_sc_hd__a22oi_1 U608 ( .A1(n10), .A2(pcgen_btb_ifpc[12]), .B1(
        pcgen_pred_ifpc[12]), .B2(n89), .Y(n387) );
  sky130_fd_sc_hd__o21ai_1 U609 ( .A1(n99), .A2(n388), .B1(n387), .Y(n445) );
  sky130_fd_sc_hd__a22oi_1 U610 ( .A1(n91), .A2(pcgen_btb_ifpc[13]), .B1(
        pcgen_pred_ifpc[13]), .B2(n90), .Y(n389) );
  sky130_fd_sc_hd__o21ai_1 U611 ( .A1(n99), .A2(n390), .B1(n389), .Y(n446) );
  sky130_fd_sc_hd__a22oi_1 U612 ( .A1(n91), .A2(pcgen_btb_ifpc[14]), .B1(
        pcgen_pred_ifpc[14]), .B2(n89), .Y(n391) );
  sky130_fd_sc_hd__o21ai_1 U613 ( .A1(n99), .A2(n392), .B1(n391), .Y(n447) );
  sky130_fd_sc_hd__a22oi_1 U614 ( .A1(n91), .A2(pcgen_btb_ifpc[15]), .B1(
        pcgen_pred_ifpc[15]), .B2(n90), .Y(n393) );
  sky130_fd_sc_hd__o21ai_1 U615 ( .A1(n99), .A2(n394), .B1(n393), .Y(n448) );
  sky130_fd_sc_hd__a22oi_1 U616 ( .A1(n91), .A2(pcgen_icache_va[16]), .B1(
        pcgen_pred_ifpc[16]), .B2(n90), .Y(n395) );
  sky130_fd_sc_hd__o21ai_1 U617 ( .A1(n99), .A2(n396), .B1(n395), .Y(n449) );
  sky130_fd_sc_hd__a22oi_1 U618 ( .A1(n91), .A2(pcgen_icache_va[17]), .B1(
        pcgen_pred_ifpc[17]), .B2(n89), .Y(n397) );
  sky130_fd_sc_hd__o21ai_1 U619 ( .A1(n98), .A2(n398), .B1(n397), .Y(n450) );
  sky130_fd_sc_hd__a22oi_1 U620 ( .A1(n91), .A2(pcgen_icache_va[18]), .B1(
        pcgen_pred_ifpc[18]), .B2(n90), .Y(n399) );
  sky130_fd_sc_hd__o21ai_1 U621 ( .A1(n98), .A2(n400), .B1(n399), .Y(n451) );
  sky130_fd_sc_hd__a22oi_1 U622 ( .A1(n10), .A2(pcgen_icache_va[19]), .B1(
        pcgen_pred_ifpc[19]), .B2(n27), .Y(n401) );
  sky130_fd_sc_hd__o21ai_1 U623 ( .A1(n98), .A2(n402), .B1(n401), .Y(n452) );
  sky130_fd_sc_hd__a22oi_1 U624 ( .A1(n91), .A2(pcgen_icache_va[20]), .B1(
        pcgen_pred_ifpc[20]), .B2(n90), .Y(n403) );
  sky130_fd_sc_hd__o21ai_1 U625 ( .A1(n98), .A2(n404), .B1(n403), .Y(n453) );
  sky130_fd_sc_hd__a22oi_1 U626 ( .A1(n91), .A2(pcgen_icache_va[21]), .B1(
        pcgen_pred_ifpc[21]), .B2(n89), .Y(n405) );
  sky130_fd_sc_hd__o21ai_1 U627 ( .A1(n98), .A2(n406), .B1(n405), .Y(n454) );
  sky130_fd_sc_hd__a22oi_1 U628 ( .A1(n10), .A2(pcgen_icache_va[22]), .B1(
        pcgen_pred_ifpc[22]), .B2(n89), .Y(n407) );
  sky130_fd_sc_hd__o21ai_1 U629 ( .A1(n98), .A2(n408), .B1(n407), .Y(n455) );
  sky130_fd_sc_hd__a22oi_1 U630 ( .A1(n92), .A2(pcgen_icache_va[23]), .B1(
        pcgen_pred_ifpc[23]), .B2(n27), .Y(n409) );
  sky130_fd_sc_hd__o21ai_1 U631 ( .A1(n99), .A2(n410), .B1(n409), .Y(n456) );
  sky130_fd_sc_hd__a22oi_1 U632 ( .A1(n93), .A2(pcgen_icache_va[24]), .B1(
        pcgen_pred_ifpc[24]), .B2(n90), .Y(n411) );
  sky130_fd_sc_hd__o21ai_1 U633 ( .A1(n99), .A2(n412), .B1(n411), .Y(n457) );
  sky130_fd_sc_hd__a22oi_1 U634 ( .A1(n11), .A2(pcgen_icache_va[25]), .B1(
        pcgen_pred_ifpc[25]), .B2(n89), .Y(n413) );
  sky130_fd_sc_hd__o21ai_1 U635 ( .A1(n98), .A2(n414), .B1(n413), .Y(n458) );
  sky130_fd_sc_hd__a22oi_1 U636 ( .A1(n92), .A2(pcgen_icache_va[26]), .B1(
        pcgen_pred_ifpc[26]), .B2(n88), .Y(n415) );
  sky130_fd_sc_hd__o21ai_1 U637 ( .A1(n98), .A2(n416), .B1(n415), .Y(n459) );
  sky130_fd_sc_hd__a22oi_1 U638 ( .A1(n93), .A2(pcgen_icache_va[27]), .B1(
        pcgen_pred_ifpc[27]), .B2(n88), .Y(n417) );
  sky130_fd_sc_hd__o21ai_1 U639 ( .A1(n98), .A2(n418), .B1(n417), .Y(n460) );
  sky130_fd_sc_hd__a22oi_1 U640 ( .A1(n11), .A2(pcgen_icache_va[28]), .B1(
        pcgen_pred_ifpc[28]), .B2(n88), .Y(n419) );
  sky130_fd_sc_hd__o21ai_1 U641 ( .A1(n98), .A2(n420), .B1(n419), .Y(n461) );
  sky130_fd_sc_hd__a22oi_1 U642 ( .A1(n10), .A2(pcgen_icache_va[29]), .B1(
        pcgen_pred_ifpc[29]), .B2(n88), .Y(n421) );
  sky130_fd_sc_hd__o21ai_1 U643 ( .A1(n98), .A2(n422), .B1(n421), .Y(n462) );
  sky130_fd_sc_hd__a22oi_1 U644 ( .A1(n92), .A2(pcgen_icache_va[30]), .B1(
        pcgen_pred_ifpc[30]), .B2(n88), .Y(n423) );
  sky130_fd_sc_hd__o21ai_1 U645 ( .A1(n98), .A2(n424), .B1(n423), .Y(n463) );
  sky130_fd_sc_hd__a22oi_1 U646 ( .A1(n93), .A2(pcgen_icache_va[31]), .B1(
        pcgen_pred_ifpc[31]), .B2(n88), .Y(n425) );
  sky130_fd_sc_hd__o21ai_1 U647 ( .A1(n98), .A2(n426), .B1(n425), .Y(n464) );
  sky130_fd_sc_hd__a22oi_1 U648 ( .A1(n11), .A2(pcgen_icache_va[32]), .B1(
        pcgen_pred_ifpc[32]), .B2(n88), .Y(n427) );
  sky130_fd_sc_hd__o21ai_1 U649 ( .A1(n98), .A2(n428), .B1(n427), .Y(n465) );
  sky130_fd_sc_hd__a22oi_1 U650 ( .A1(n92), .A2(pcgen_icache_va[33]), .B1(
        pcgen_pred_ifpc[33]), .B2(n90), .Y(n429) );
  sky130_fd_sc_hd__o21ai_1 U651 ( .A1(n99), .A2(n430), .B1(n429), .Y(n466) );
  sky130_fd_sc_hd__a22oi_1 U652 ( .A1(n92), .A2(pcgen_icache_va[34]), .B1(
        pcgen_pred_ifpc[34]), .B2(n90), .Y(n431) );
  sky130_fd_sc_hd__o21ai_1 U653 ( .A1(n98), .A2(n432), .B1(n431), .Y(n467) );
  sky130_fd_sc_hd__a22oi_1 U654 ( .A1(n93), .A2(pcgen_icache_va[35]), .B1(
        pcgen_pred_ifpc[35]), .B2(n89), .Y(n473) );
  sky130_fd_sc_hd__o21ai_1 U655 ( .A1(n98), .A2(n474), .B1(n473), .Y(n468) );
  sky130_fd_sc_hd__a22oi_1 U656 ( .A1(n11), .A2(pcgen_icache_va[36]), .B1(
        pcgen_pred_ifpc[36]), .B2(n88), .Y(n475) );
  sky130_fd_sc_hd__o21ai_1 U657 ( .A1(n98), .A2(n476), .B1(n475), .Y(n469) );
  sky130_fd_sc_hd__a22oi_1 U658 ( .A1(n10), .A2(pcgen_icache_va[37]), .B1(
        pcgen_pred_ifpc[37]), .B2(n27), .Y(n477) );
  sky130_fd_sc_hd__o21ai_1 U659 ( .A1(n99), .A2(n478), .B1(n477), .Y(n470) );
  sky130_fd_sc_hd__a22oi_1 U660 ( .A1(n93), .A2(pcgen_icache_va[38]), .B1(
        pcgen_pred_ifpc[38]), .B2(n89), .Y(n481) );
  sky130_fd_sc_hd__o21ai_1 U661 ( .A1(n98), .A2(n482), .B1(n481), .Y(n471) );
  sky130_fd_sc_hd__inv_1 U662 ( .A(pcgen_pred_ifpc[39]), .Y(n484) );
  sky130_fd_sc_hd__o221ai_1 U663 ( .A1(n487), .A2(n9), .B1(n8), .B2(n484), 
        .C1(n483), .Y(n472) );
  sky130_fd_sc_hd__inv_1 U664 ( .A(btb_xx_chgflw_vld), .Y(n489) );
  sky130_fd_sc_hd__nand3_1 U665 ( .A(n28), .B(n489), .C(n55), .Y(
        pcgen_icache_chgflw_vld) );
endmodule


module aq_ifu_ctrl_0 ( cp0_ifu_in_lpmd, cp0_ifu_lpmd_req, ctrl_btb_chgflw_vld, 
        ctrl_btb_inst_fetch, ctrl_btb_stall, ctrl_ibuf_pop_en, 
        ctrl_icache_abort, ctrl_icache_req_vld, ctrl_ipack_cancel, 
        ibuf_ctrl_inst_fetch, icache_ctrl_stall, idu_ifu_id_stall, 
        pcgen_ctrl_chgflw_vld, pred_ctrl_stall, rtu_ifu_dbg_mask, 
        rtu_ifu_flush_fe, vec_ctrl_reset_mask );
  input cp0_ifu_in_lpmd, cp0_ifu_lpmd_req, ibuf_ctrl_inst_fetch,
         icache_ctrl_stall, idu_ifu_id_stall, pcgen_ctrl_chgflw_vld,
         pred_ctrl_stall, rtu_ifu_dbg_mask, rtu_ifu_flush_fe,
         vec_ctrl_reset_mask;
  output ctrl_btb_chgflw_vld, ctrl_btb_inst_fetch, ctrl_btb_stall,
         ctrl_ibuf_pop_en, ctrl_icache_abort, ctrl_icache_req_vld,
         ctrl_ipack_cancel;
  wire   ctrl_icache_abort, ctrl_icache_req_vld, n3;
  assign ctrl_btb_chgflw_vld = ctrl_icache_abort;
  assign ctrl_btb_inst_fetch = ctrl_icache_req_vld;

  sky130_fd_sc_hd__nor4_4 U1 ( .A(rtu_ifu_dbg_mask), .B(n3), .C(
        cp0_ifu_in_lpmd), .D(cp0_ifu_lpmd_req), .Y(ctrl_icache_req_vld) );
  sky130_fd_sc_hd__or2_4 U2 ( .A(rtu_ifu_flush_fe), .B(pcgen_ctrl_chgflw_vld), 
        .X(ctrl_icache_abort) );
  sky130_fd_sc_hd__or2_1 U3 ( .A(rtu_ifu_flush_fe), .B(pcgen_ctrl_chgflw_vld), 
        .X(ctrl_ipack_cancel) );
  sky130_fd_sc_hd__nand2b_1 U4 ( .A_N(vec_ctrl_reset_mask), .B(
        ibuf_ctrl_inst_fetch), .Y(n3) );
  sky130_fd_sc_hd__inv_1 U5 ( .A(idu_ifu_id_stall), .Y(ctrl_ibuf_pop_en) );
  sky130_fd_sc_hd__or2_0 U6 ( .A(icache_ctrl_stall), .B(pred_ctrl_stall), .X(
        ctrl_btb_stall) );
endmodule