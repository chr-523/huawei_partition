
module aq_iu_mul_0_DW01_add_5 ( A, B, CI, SUM, CO );
  input [68:0] A;
  input [68:0] B;
  output [68:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n8, n13, n14, n15, n16, n17, n18, n19, n20, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201;
  assign SUM[0] = B[0];

  sky130_fd_sc_hd__inv_1 U2 ( .A(n62), .Y(n84) );
  sky130_fd_sc_hd__clkinv_1 U3 ( .A(n81), .Y(n74) );
  sky130_fd_sc_hd__inv_1 U4 ( .A(n131), .Y(n144) );
  sky130_fd_sc_hd__clkinv_1 U5 ( .A(n73), .Y(n72) );
  sky130_fd_sc_hd__inv_1 U6 ( .A(n200), .Y(n36) );
  sky130_fd_sc_hd__inv_1 U7 ( .A(n195), .Y(n53) );
  sky130_fd_sc_hd__inv_1 U8 ( .A(n143), .Y(n141) );
  sky130_fd_sc_hd__inv_1 U9 ( .A(n71), .Y(n68) );
  sky130_fd_sc_hd__inv_1 U10 ( .A(n113), .Y(n112) );
  sky130_fd_sc_hd__xor2_2 U11 ( .A(n57), .B(B[67]), .X(SUM[67]) );
  sky130_fd_sc_hd__clkinv_1 U12 ( .A(n162), .Y(n154) );
  sky130_fd_sc_hd__inv_2 U13 ( .A(n75), .Y(n48) );
  sky130_fd_sc_hd__and2_1 U14 ( .A(B[30]), .B(B[28]), .X(n135) );
  sky130_fd_sc_hd__inv_1 U15 ( .A(B[20]), .Y(n153) );
  sky130_fd_sc_hd__and2_1 U16 ( .A(n8), .B(B[49]), .X(n20) );
  sky130_fd_sc_hd__and2_1 U17 ( .A(B[1]), .B(A[1]), .X(n34) );
  sky130_fd_sc_hd__inv_1 U18 ( .A(n128), .Y(n90) );
  sky130_fd_sc_hd__inv_1 U19 ( .A(n44), .Y(n117) );
  sky130_fd_sc_hd__inv_1 U20 ( .A(n169), .Y(n162) );
  sky130_fd_sc_hd__inv_1 U21 ( .A(n109), .Y(n108) );
  sky130_fd_sc_hd__and2_1 U22 ( .A(n144), .B(n145), .X(n5) );
  sky130_fd_sc_hd__clkinv_1 U23 ( .A(n163), .Y(n150) );
  sky130_fd_sc_hd__inv_1 U24 ( .A(n95), .Y(n124) );
  sky130_fd_sc_hd__inv_1 U25 ( .A(n161), .Y(n156) );
  sky130_fd_sc_hd__and2_1 U26 ( .A(n5), .B(B[28]), .X(n13) );
  sky130_fd_sc_hd__and2_1 U27 ( .A(n19), .B(n68), .X(n18) );
  sky130_fd_sc_hd__and2_1 U28 ( .A(B[57]), .B(n15), .X(n80) );
  sky130_fd_sc_hd__and2_1 U29 ( .A(B[53]), .B(n16), .X(n83) );
  sky130_fd_sc_hd__inv_1 U30 ( .A(n132), .Y(n151) );
  sky130_fd_sc_hd__and2_1 U31 ( .A(n3), .B(B[64]), .X(n14) );
  sky130_fd_sc_hd__and2_1 U32 ( .A(n17), .B(B[52]), .X(n16) );
  sky130_fd_sc_hd__and2_1 U33 ( .A(B[65]), .B(n14), .X(n58) );
  sky130_fd_sc_hd__and2_1 U34 ( .A(n74), .B(B[56]), .X(n15) );
  sky130_fd_sc_hd__and2_1 U35 ( .A(n72), .B(B[60]), .X(n19) );
  sky130_fd_sc_hd__inv_1 U36 ( .A(n191), .Y(n183) );
  sky130_fd_sc_hd__inv_1 U37 ( .A(n39), .Y(n191) );
  sky130_fd_sc_hd__clkinv_1 U38 ( .A(n78), .Y(n77) );
  sky130_fd_sc_hd__xor2_1 U39 ( .A(n1), .B(B[23]), .X(SUM[23]) );
  sky130_fd_sc_hd__nor2_1 U40 ( .A(n154), .B(n155), .Y(n1) );
  sky130_fd_sc_hd__xor2_1 U41 ( .A(n2), .B(B[21]), .X(SUM[21]) );
  sky130_fd_sc_hd__nor2_1 U42 ( .A(n169), .B(n161), .Y(n2) );
  sky130_fd_sc_hd__and2_1 U43 ( .A(n111), .B(B[41]), .X(n28) );
  sky130_fd_sc_hd__and2_1 U44 ( .A(n30), .B(B[37]), .X(n29) );
  sky130_fd_sc_hd__and2_1 U45 ( .A(B[33]), .B(n127), .X(n126) );
  sky130_fd_sc_hd__and2_1 U46 ( .A(B[48]), .B(n60), .X(n8) );
  sky130_fd_sc_hd__and2_1 U47 ( .A(B[36]), .B(n114), .X(n30) );
  sky130_fd_sc_hd__and2_1 U48 ( .A(n142), .B(n178), .X(SUM[1]) );
  sky130_fd_sc_hd__xnor2_1 U49 ( .A(n186), .B(B[13]), .Y(SUM[13]) );
  sky130_fd_sc_hd__xor2_1 U50 ( .A(n200), .B(n39), .X(SUM[8]) );
  sky130_fd_sc_hd__xor2_1 U51 ( .A(n35), .B(n201), .X(SUM[9]) );
  sky130_fd_sc_hd__xor2_1 U52 ( .A(n197), .B(n196), .X(SUM[10]) );
  sky130_fd_sc_hd__inv_1 U53 ( .A(B[12]), .Y(n189) );
  sky130_fd_sc_hd__xor2_1 U54 ( .A(n78), .B(n46), .X(SUM[4]) );
  sky130_fd_sc_hd__inv_1 U55 ( .A(n176), .Y(n184) );
  sky130_fd_sc_hd__inv_1 U56 ( .A(B[14]), .Y(n180) );
  sky130_fd_sc_hd__inv_1 U57 ( .A(B[45]), .Y(n100) );
  sky130_fd_sc_hd__inv_1 U58 ( .A(B[44]), .Y(n98) );
  sky130_fd_sc_hd__inv_1 U59 ( .A(n177), .Y(n176) );
  sky130_fd_sc_hd__inv_1 U60 ( .A(n38), .Y(n37) );
  sky130_fd_sc_hd__inv_1 U61 ( .A(n55), .Y(n49) );
  sky130_fd_sc_hd__xor2_1 U62 ( .A(n181), .B(n180), .X(SUM[14]) );
  sky130_fd_sc_hd__nor2_1 U63 ( .A(n90), .B(n91), .Y(n60) );
  sky130_fd_sc_hd__nor2_1 U64 ( .A(n101), .B(n102), .Y(n92) );
  sky130_fd_sc_hd__nor2_1 U65 ( .A(n113), .B(n101), .Y(n109) );
  sky130_fd_sc_hd__nor2_1 U66 ( .A(n169), .B(n122), .Y(n128) );
  sky130_fd_sc_hd__nor2_1 U67 ( .A(n90), .B(n99), .Y(n127) );
  sky130_fd_sc_hd__nor2_1 U68 ( .A(n98), .B(n108), .Y(n107) );
  sky130_fd_sc_hd__nor2_1 U69 ( .A(n143), .B(n140), .Y(n139) );
  sky130_fd_sc_hd__inv_2 U70 ( .A(n13), .Y(n140) );
  sky130_fd_sc_hd__nor2_1 U71 ( .A(n100), .B(n106), .Y(n105) );
  sky130_fd_sc_hd__inv_1 U72 ( .A(n107), .Y(n106) );
  sky130_fd_sc_hd__nor2_1 U73 ( .A(n169), .B(n147), .Y(n145) );
  sky130_fd_sc_hd__nor2_1 U74 ( .A(n180), .B(n181), .Y(n179) );
  sky130_fd_sc_hd__nor3_1 U75 ( .A(n62), .B(n63), .C(n64), .Y(n61) );
  sky130_fd_sc_hd__nand2b_1 U76 ( .A_N(n102), .B(n114), .Y(n113) );
  sky130_fd_sc_hd__nand2b_1 U77 ( .A_N(n64), .B(n17), .Y(n81) );
  sky130_fd_sc_hd__nor2_1 U78 ( .A(n4), .B(n59), .Y(n3) );
  sky130_fd_sc_hd__or2_2 U79 ( .A(n65), .B(n66), .X(n4) );
  sky130_fd_sc_hd__nand2b_1 U80 ( .A_N(n63), .B(n74), .Y(n73) );
  sky130_fd_sc_hd__xnor2_1 U81 ( .A(n190), .B(n189), .Y(SUM[12]) );
  sky130_fd_sc_hd__nor2_1 U82 ( .A(n183), .B(n184), .Y(n190) );
  sky130_fd_sc_hd__xnor2_1 U83 ( .A(n164), .B(n153), .Y(SUM[20]) );
  sky130_fd_sc_hd__nor2_1 U84 ( .A(n169), .B(n163), .Y(n164) );
  sky130_fd_sc_hd__xor2_1 U85 ( .A(n116), .B(n117), .X(SUM[2]) );
  sky130_fd_sc_hd__nor2_1 U86 ( .A(n189), .B(n184), .Y(n187) );
  sky130_fd_sc_hd__xor2_1 U87 ( .A(n103), .B(n104), .X(SUM[47]) );
  sky130_fd_sc_hd__xor2_1 U88 ( .A(n80), .B(B[58]), .X(SUM[58]) );
  sky130_fd_sc_hd__xor2_1 U89 ( .A(n137), .B(n138), .X(SUM[31]) );
  sky130_fd_sc_hd__xnor2_1 U90 ( .A(n159), .B(n158), .Y(SUM[22]) );
  sky130_fd_sc_hd__nor2_1 U91 ( .A(n154), .B(n160), .Y(n159) );
  sky130_fd_sc_hd__xor2_1 U92 ( .A(n83), .B(B[54]), .X(SUM[54]) );
  sky130_fd_sc_hd__xor2_1 U93 ( .A(n105), .B(B[46]), .X(SUM[46]) );
  sky130_fd_sc_hd__xnor2_1 U94 ( .A(n76), .B(n48), .Y(SUM[5]) );
  sky130_fd_sc_hd__xor2_1 U95 ( .A(n58), .B(B[66]), .X(SUM[66]) );
  sky130_fd_sc_hd__xor2_1 U96 ( .A(n69), .B(n70), .X(SUM[63]) );
  sky130_fd_sc_hd__xor2_1 U97 ( .A(n13), .B(n141), .X(SUM[29]) );
  sky130_fd_sc_hd__xor2_1 U98 ( .A(n15), .B(B[57]), .X(SUM[57]) );
  sky130_fd_sc_hd__xor2_1 U99 ( .A(n14), .B(B[65]), .X(SUM[65]) );
  sky130_fd_sc_hd__xor2_1 U100 ( .A(n74), .B(B[56]), .X(SUM[56]) );
  sky130_fd_sc_hd__xor2_1 U101 ( .A(n3), .B(B[64]), .X(SUM[64]) );
  sky130_fd_sc_hd__xor2_1 U102 ( .A(n18), .B(B[62]), .X(SUM[62]) );
  sky130_fd_sc_hd__xor2_1 U103 ( .A(n139), .B(B[30]), .X(SUM[30]) );
  sky130_fd_sc_hd__xor2_1 U104 ( .A(n19), .B(n68), .X(SUM[61]) );
  sky130_fd_sc_hd__xor2_1 U105 ( .A(n5), .B(B[28]), .X(SUM[28]) );
  sky130_fd_sc_hd__xor2_1 U106 ( .A(n20), .B(B[50]), .X(SUM[50]) );
  sky130_fd_sc_hd__xor2_1 U107 ( .A(n126), .B(B[34]), .X(SUM[34]) );
  sky130_fd_sc_hd__xnor2_1 U108 ( .A(B[55]), .B(n82), .Y(SUM[55]) );
  sky130_fd_sc_hd__and2_0 U109 ( .A(B[66]), .B(n58), .X(n57) );
  sky130_fd_sc_hd__nand2b_1 U110 ( .A_N(n134), .B(B[16]), .Y(n163) );
  sky130_fd_sc_hd__nor2_1 U111 ( .A(n169), .B(n167), .Y(n166) );
  sky130_fd_sc_hd__nor2_1 U112 ( .A(n184), .B(n185), .Y(n182) );
  sky130_fd_sc_hd__nor2_1 U113 ( .A(n131), .B(n132), .Y(n130) );
  sky130_fd_sc_hd__nand3_1 U114 ( .A(n135), .B(n136), .C(B[16]), .Y(n133) );
  sky130_fd_sc_hd__nor2_1 U115 ( .A(n138), .B(n143), .Y(n136) );
  sky130_fd_sc_hd__xnor2_1 U116 ( .A(B[59]), .B(n79), .Y(SUM[59]) );
  sky130_fd_sc_hd__nand3_1 U117 ( .A(B[17]), .B(B[19]), .C(B[18]), .Y(n134) );
  sky130_fd_sc_hd__nand3_1 U118 ( .A(B[33]), .B(B[35]), .C(B[34]), .Y(n95) );
  sky130_fd_sc_hd__clkinv_1 U119 ( .A(n169), .Y(n120) );
  sky130_fd_sc_hd__nor2_1 U120 ( .A(n172), .B(n173), .Y(n171) );
  sky130_fd_sc_hd__nor2_1 U121 ( .A(n174), .B(n175), .Y(n170) );
  sky130_fd_sc_hd__xor2_1 U122 ( .A(B[15]), .B(n179), .X(SUM[15]) );
  sky130_fd_sc_hd__xnor2_1 U123 ( .A(B[19]), .B(n165), .Y(SUM[19]) );
  sky130_fd_sc_hd__xnor2_1 U124 ( .A(B[35]), .B(n125), .Y(SUM[35]) );
  sky130_fd_sc_hd__xnor2_1 U125 ( .A(B[51]), .B(n85), .Y(SUM[51]) );
  sky130_fd_sc_hd__clkinv_1 U126 ( .A(n119), .Y(n114) );
  sky130_fd_sc_hd__nor2_1 U127 ( .A(n122), .B(n123), .Y(n121) );
  sky130_fd_sc_hd__and3_1 U128 ( .A(B[48]), .B(n84), .C(n60), .X(n17) );
  sky130_fd_sc_hd__xor2_1 U129 ( .A(n72), .B(B[60]), .X(SUM[60]) );
  sky130_fd_sc_hd__xor2_1 U130 ( .A(n16), .B(B[53]), .X(SUM[53]) );
  sky130_fd_sc_hd__xor2_1 U131 ( .A(n107), .B(B[45]), .X(SUM[45]) );
  sky130_fd_sc_hd__xor2_1 U132 ( .A(n127), .B(B[33]), .X(SUM[33]) );
  sky130_fd_sc_hd__xor2_1 U133 ( .A(n8), .B(B[49]), .X(SUM[49]) );
  sky130_fd_sc_hd__xor2_1 U134 ( .A(n30), .B(B[37]), .X(SUM[37]) );
  sky130_fd_sc_hd__xor2_1 U135 ( .A(n166), .B(B[18]), .X(SUM[18]) );
  sky130_fd_sc_hd__xor2_1 U136 ( .A(n27), .B(B[26]), .X(SUM[26]) );
  sky130_fd_sc_hd__xor2_1 U137 ( .A(n109), .B(B[44]), .X(SUM[44]) );
  sky130_fd_sc_hd__xor2_1 U138 ( .A(n145), .B(B[24]), .X(SUM[24]) );
  sky130_fd_sc_hd__xor2_1 U139 ( .A(n17), .B(B[52]), .X(SUM[52]) );
  sky130_fd_sc_hd__xor2_1 U140 ( .A(n60), .B(B[48]), .X(SUM[48]) );
  sky130_fd_sc_hd__xor2_1 U141 ( .A(n112), .B(B[40]), .X(SUM[40]) );
  sky130_fd_sc_hd__xor2_1 U142 ( .A(n120), .B(B[16]), .X(SUM[16]) );
  sky130_fd_sc_hd__xor2_1 U143 ( .A(n128), .B(B[32]), .X(SUM[32]) );
  sky130_fd_sc_hd__xor2_1 U144 ( .A(n114), .B(B[36]), .X(SUM[36]) );
  sky130_fd_sc_hd__xor2_1 U145 ( .A(n28), .B(B[42]), .X(SUM[42]) );
  sky130_fd_sc_hd__xor2_1 U146 ( .A(n29), .B(B[38]), .X(SUM[38]) );
  sky130_fd_sc_hd__xor2_1 U147 ( .A(n111), .B(B[41]), .X(SUM[41]) );
  sky130_fd_sc_hd__nor2b_1 U148 ( .B_N(B[40]), .A(n113), .Y(n111) );
  sky130_fd_sc_hd__nor3_1 U149 ( .A(n195), .B(n196), .C(n44), .Y(n194) );
  sky130_fd_sc_hd__nor2b_1 U150 ( .B_N(n49), .A(n195), .Y(n41) );
  sky130_fd_sc_hd__nand3_1 U151 ( .A(B[49]), .B(B[51]), .C(B[50]), .Y(n62) );
  sky130_fd_sc_hd__nand3_1 U152 ( .A(B[24]), .B(n149), .C(n120), .Y(n148) );
  sky130_fd_sc_hd__inv_1 U153 ( .A(n147), .Y(n149) );
  sky130_fd_sc_hd__nor2b_1 U154 ( .B_N(B[21]), .A(n158), .Y(n157) );
  sky130_fd_sc_hd__nor2_1 U155 ( .A(n200), .B(n201), .Y(n193) );
  sky130_fd_sc_hd__xnor2_1 U156 ( .A(B[27]), .B(n146), .Y(SUM[27]) );
  sky130_fd_sc_hd__xnor2_1 U157 ( .A(B[43]), .B(n110), .Y(SUM[43]) );
  sky130_fd_sc_hd__xnor2_1 U158 ( .A(B[39]), .B(n118), .Y(SUM[39]) );
  sky130_fd_sc_hd__xor2_1 U159 ( .A(n49), .B(n50), .X(SUM[6]) );
  sky130_fd_sc_hd__xnor2_1 U160 ( .A(n148), .B(B[25]), .Y(SUM[25]) );
  sky130_fd_sc_hd__xnor2_1 U161 ( .A(n168), .B(B[17]), .Y(SUM[17]) );
  sky130_fd_sc_hd__inv_1 U162 ( .A(n142), .Y(n116) );
  sky130_fd_sc_hd__nand3_1 U163 ( .A(n96), .B(B[46]), .C(n97), .Y(n94) );
  sky130_fd_sc_hd__nor2_1 U164 ( .A(n104), .B(n100), .Y(n96) );
  sky130_fd_sc_hd__nor2_1 U165 ( .A(n98), .B(n99), .Y(n97) );
  sky130_fd_sc_hd__inv_2 U166 ( .A(n54), .Y(n46) );
  sky130_fd_sc_hd__and4_1 U167 ( .A(B[24]), .B(B[25]), .C(n149), .D(n120), .X(
        n27) );
  sky130_fd_sc_hd__nor2_1 U168 ( .A(n70), .B(n71), .Y(n67) );
  sky130_fd_sc_hd__inv_2 U169 ( .A(B[32]), .Y(n99) );
  sky130_fd_sc_hd__inv_1 U170 ( .A(n39), .Y(n188) );
  sky130_fd_sc_hd__inv_2 U171 ( .A(n48), .Y(n47) );
  sky130_fd_sc_hd__and4_1 U172 ( .A(B[3]), .B(B[1]), .C(A[1]), .D(B[2]), .X(
        n31) );
  sky130_fd_sc_hd__and4_1 U173 ( .A(B[7]), .B(B[6]), .C(B[5]), .D(B[4]), .X(
        n32) );
  sky130_fd_sc_hd__nand3_1 U174 ( .A(B[2]), .B(n53), .C(n87), .Y(n78) );
  sky130_fd_sc_hd__inv_1 U175 ( .A(B[2]), .Y(n44) );
  sky130_fd_sc_hd__nand3_1 U176 ( .A(B[1]), .B(A[1]), .C(B[3]), .Y(n198) );
  sky130_fd_sc_hd__nor3_1 U177 ( .A(n44), .B(n201), .C(n200), .Y(n199) );
  sky130_fd_sc_hd__nand3_1 U178 ( .A(B[23]), .B(n152), .C(B[21]), .Y(n132) );
  sky130_fd_sc_hd__nor2_1 U179 ( .A(n153), .B(n158), .Y(n152) );
  sky130_fd_sc_hd__inv_1 U180 ( .A(A[1]), .Y(n88) );
  sky130_fd_sc_hd__inv_1 U181 ( .A(B[1]), .Y(n89) );
  sky130_fd_sc_hd__nand3_1 U182 ( .A(B[4]), .B(B[6]), .C(B[5]), .Y(n173) );
  sky130_fd_sc_hd__inv_1 U183 ( .A(B[22]), .Y(n158) );
  sky130_fd_sc_hd__inv_1 U184 ( .A(B[3]), .Y(n195) );
  sky130_fd_sc_hd__inv_1 U185 ( .A(B[31]), .Y(n138) );
  sky130_fd_sc_hd__inv_1 U186 ( .A(B[29]), .Y(n143) );
  sky130_fd_sc_hd__xnor2_1 U187 ( .A(n192), .B(B[11]), .Y(SUM[11]) );
  sky130_fd_sc_hd__xor2_1 U188 ( .A(n115), .B(n195), .X(SUM[3]) );
  sky130_fd_sc_hd__nand3_1 U189 ( .A(n41), .B(n42), .C(n43), .Y(n40) );
  sky130_fd_sc_hd__nor2_1 U190 ( .A(n46), .B(n47), .Y(n42) );
  sky130_fd_sc_hd__nor2_1 U191 ( .A(n51), .B(n52), .Y(n50) );
  sky130_fd_sc_hd__and4_1 U192 ( .A(B[7]), .B(B[6]), .C(B[5]), .D(B[4]), .X(
        n33) );
  sky130_fd_sc_hd__inv_1 U193 ( .A(B[5]), .Y(n75) );
  sky130_fd_sc_hd__inv_1 U194 ( .A(B[6]), .Y(n55) );
  sky130_fd_sc_hd__inv_2 U195 ( .A(n86), .Y(n54) );
  sky130_fd_sc_hd__inv_1 U196 ( .A(B[4]), .Y(n86) );
  sky130_fd_sc_hd__inv_1 U197 ( .A(B[63]), .Y(n70) );
  sky130_fd_sc_hd__inv_1 U198 ( .A(B[47]), .Y(n104) );
  sky130_fd_sc_hd__inv_1 U199 ( .A(B[10]), .Y(n196) );
  sky130_fd_sc_hd__inv_1 U200 ( .A(B[9]), .Y(n201) );
  sky130_fd_sc_hd__inv_1 U201 ( .A(B[8]), .Y(n200) );
  sky130_fd_sc_hd__inv_1 U202 ( .A(B[61]), .Y(n71) );
  sky130_fd_sc_hd__nand2_1 U203 ( .A(n116), .B(n117), .Y(n115) );
  sky130_fd_sc_hd__nand2_1 U204 ( .A(n57), .B(B[67]), .Y(n56) );
  sky130_fd_sc_hd__nand2_1 U205 ( .A(n18), .B(B[62]), .Y(n69) );
  sky130_fd_sc_hd__nand2_1 U206 ( .A(n105), .B(B[46]), .Y(n103) );
  sky130_fd_sc_hd__nand2_1 U207 ( .A(n139), .B(B[30]), .Y(n137) );
  sky130_fd_sc_hd__nand2_1 U208 ( .A(n170), .B(n171), .Y(n169) );
  sky130_fd_sc_hd__nand2_1 U209 ( .A(n80), .B(B[58]), .Y(n79) );
  sky130_fd_sc_hd__nand2_1 U210 ( .A(n83), .B(B[54]), .Y(n82) );
  sky130_fd_sc_hd__nand2_1 U211 ( .A(n20), .B(B[50]), .Y(n85) );
  sky130_fd_sc_hd__nand2_1 U212 ( .A(n28), .B(B[42]), .Y(n110) );
  sky130_fd_sc_hd__nand2_1 U213 ( .A(n29), .B(B[38]), .Y(n118) );
  sky130_fd_sc_hd__nand2_1 U214 ( .A(n126), .B(B[34]), .Y(n125) );
  sky130_fd_sc_hd__nand2_1 U215 ( .A(n27), .B(B[26]), .Y(n146) );
  sky130_fd_sc_hd__nand2_1 U216 ( .A(n166), .B(B[18]), .Y(n165) );
  sky130_fd_sc_hd__nand2_1 U217 ( .A(n182), .B(n191), .Y(n181) );
  sky130_fd_sc_hd__nand2_1 U218 ( .A(n187), .B(n188), .Y(n186) );
  sky130_fd_sc_hd__nand3_1 U219 ( .A(n33), .B(n36), .C(n37), .Y(n35) );
  sky130_fd_sc_hd__nand4_1 U220 ( .A(B[3]), .B(B[1]), .C(A[1]), .D(B[2]), .Y(
        n38) );
  sky130_fd_sc_hd__xnor2_1 U221 ( .A(n40), .B(B[7]), .Y(SUM[7]) );
  sky130_fd_sc_hd__nor2_1 U222 ( .A(n44), .B(n45), .Y(n43) );
  sky130_fd_sc_hd__nand2_1 U223 ( .A(A[1]), .B(B[1]), .Y(n45) );
  sky130_fd_sc_hd__nand4_1 U224 ( .A(A[1]), .B(B[1]), .C(B[2]), .D(n53), .Y(
        n52) );
  sky130_fd_sc_hd__nand2_1 U225 ( .A(n48), .B(n54), .Y(n51) );
  sky130_fd_sc_hd__xnor2_1 U226 ( .A(n56), .B(B[68]), .Y(SUM[68]) );
  sky130_fd_sc_hd__nand2_1 U227 ( .A(n60), .B(n61), .Y(n59) );
  sky130_fd_sc_hd__nand2_1 U228 ( .A(B[48]), .B(B[60]), .Y(n66) );
  sky130_fd_sc_hd__nand2_1 U229 ( .A(n67), .B(B[62]), .Y(n65) );
  sky130_fd_sc_hd__nand4_1 U230 ( .A(B[56]), .B(B[57]), .C(B[58]), .D(B[59]), 
        .Y(n63) );
  sky130_fd_sc_hd__nand2_1 U231 ( .A(n77), .B(n54), .Y(n76) );
  sky130_fd_sc_hd__nand4_1 U232 ( .A(B[52]), .B(B[53]), .C(B[54]), .D(B[55]), 
        .Y(n64) );
  sky130_fd_sc_hd__nor2_1 U233 ( .A(n88), .B(n89), .Y(n87) );
  sky130_fd_sc_hd__nand2_1 U234 ( .A(n92), .B(n93), .Y(n91) );
  sky130_fd_sc_hd__nor2_1 U235 ( .A(n94), .B(n95), .Y(n93) );
  sky130_fd_sc_hd__nand4_1 U236 ( .A(B[41]), .B(B[40]), .C(B[42]), .D(B[43]), 
        .Y(n101) );
  sky130_fd_sc_hd__nand4_1 U237 ( .A(B[36]), .B(B[37]), .C(B[38]), .D(B[39]), 
        .Y(n102) );
  sky130_fd_sc_hd__nand2_1 U238 ( .A(n120), .B(n121), .Y(n119) );
  sky130_fd_sc_hd__nand2_1 U239 ( .A(n124), .B(B[32]), .Y(n123) );
  sky130_fd_sc_hd__nand2_1 U240 ( .A(n129), .B(n130), .Y(n122) );
  sky130_fd_sc_hd__nor2_1 U241 ( .A(n133), .B(n134), .Y(n129) );
  sky130_fd_sc_hd__nand4_1 U242 ( .A(B[25]), .B(B[24]), .C(B[26]), .D(B[27]), 
        .Y(n131) );
  sky130_fd_sc_hd__nand2_1 U243 ( .A(n150), .B(n151), .Y(n147) );
  sky130_fd_sc_hd__nand2_1 U244 ( .A(n156), .B(n157), .Y(n155) );
  sky130_fd_sc_hd__nand2_1 U245 ( .A(n156), .B(B[21]), .Y(n160) );
  sky130_fd_sc_hd__nand2_1 U246 ( .A(n150), .B(B[20]), .Y(n161) );
  sky130_fd_sc_hd__nand2_1 U247 ( .A(B[1]), .B(A[1]), .Y(n142) );
  sky130_fd_sc_hd__nand2_1 U248 ( .A(B[17]), .B(B[16]), .Y(n167) );
  sky130_fd_sc_hd__nand2_1 U249 ( .A(n120), .B(B[16]), .Y(n168) );
  sky130_fd_sc_hd__nand4_1 U250 ( .A(B[12]), .B(B[14]), .C(B[13]), .D(B[15]), 
        .Y(n172) );
  sky130_fd_sc_hd__nand4_1 U251 ( .A(B[7]), .B(B[2]), .C(A[1]), .D(n176), .Y(
        n175) );
  sky130_fd_sc_hd__nand2_1 U252 ( .A(B[3]), .B(B[1]), .Y(n174) );
  sky130_fd_sc_hd__nand2_1 U253 ( .A(B[12]), .B(B[13]), .Y(n185) );
  sky130_fd_sc_hd__nand4_1 U254 ( .A(B[10]), .B(B[11]), .C(B[9]), .D(B[8]), 
        .Y(n177) );
  sky130_fd_sc_hd__nand2_1 U255 ( .A(n31), .B(n32), .Y(n39) );
  sky130_fd_sc_hd__nand4_1 U256 ( .A(n193), .B(n34), .C(n32), .D(n194), .Y(
        n192) );
  sky130_fd_sc_hd__nand3b_1 U257 ( .A_N(n198), .B(n199), .C(n32), .Y(n197) );
  sky130_fd_sc_hd__nand2_1 U258 ( .A(n89), .B(n88), .Y(n178) );
endmodule
